/*************************************************************************
   > File Name: dig_top.sv
   > Author: dafei.xiao
   > Mail: dafei.xiao@joulwatt.com
   > Created Time: Thu Sep 14 13:32:13 2023
 ************************************************************************/

module dig_top();

endmodule
