/*************************************************************************
   > File Name: adc_top.sv
   > Author: dafei.xiao
   > Mail: dafei.xiao@joulwatt.com
   > Created Time: Thu Sep 14 13:30:16 2023
 ************************************************************************/
module adc_top(






);


endmodule

