/*************************************************************************
   > File Name: system.sv
   > Author: dafei.xiao
   > Mail: dafei.xiao@joulwatt.com
   > Created Time: Thu Sep 14 13:31:34 2023
 ************************************************************************/
`include "../8_hdl/system/system.sv"

