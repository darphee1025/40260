
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.5.110
#
# REF LIBS: A11 
# TECH LIB NAME: A11
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

#NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;


PROPERTYDEFINITIONS
    LAYER LEF57_ARRAYSPACING STRING ;
    LAYER LEF57_SPACING STRING ;

END PROPERTYDEFINITIONS
 USEMINSPACING PIN OFF  ;
 USEMINSPACING OBS OFF  ;
 CLEARANCEMEASURE EUCLIDEAN  ;

SITE CORE_6T
    SYMMETRY Y    ;
    CLASS CORE  ;
    SIZE 0.400 BY 2.400 ;
END CORE_6T

SITE CORE_6T2
    SYMMETRY Y    ;
    CLASS CORE  ;
    SIZE 0.400 BY 4.800 ;
END CORE_6T2

MACRO XOR4M4HM
    CLASS CORE ;
    FOREIGN XOR4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.850 1.100 11.100 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.040 1.130 8.520 1.500 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.750 3.560 1.120 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.232  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.030 0.700 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.644  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 1.240 7.660 2.080 ;
        RECT  7.380 0.640 7.660 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  10.830 1.780 11.030 2.540 ;
        RECT  7.940 1.840 8.140 2.540 ;
        RECT  6.690 1.800 6.850 2.540 ;
        RECT  3.930 1.800 4.130 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  10.840 -0.140 11.040 0.600 ;
        RECT  8.140 -0.140 8.340 0.640 ;
        RECT  6.700 -0.140 6.900 0.570 ;
        RECT  3.400 -0.140 3.600 0.560 ;
        RECT  0.660 -0.140 0.860 0.750 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.650 1.620 1.760 ;
        RECT  1.420 1.540 1.700 1.760 ;
        RECT  0.140 0.470 0.340 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.860 1.280 2.060 2.080 ;
        RECT  1.100 1.920 2.060 2.080 ;
        RECT  1.820 0.640 1.980 1.120 ;
        RECT  1.820 0.960 2.380 1.120 ;
        RECT  2.220 0.960 2.380 2.080 ;
        RECT  2.220 1.920 2.750 2.080 ;
        RECT  1.020 0.320 3.060 0.480 ;
        RECT  2.900 0.320 3.060 1.440 ;
        RECT  1.020 0.320 1.180 1.350 ;
        RECT  2.900 1.280 3.450 1.440 ;
        RECT  3.290 1.280 3.450 1.760 ;
        RECT  2.140 0.640 2.740 0.800 ;
        RECT  2.540 0.640 2.740 1.760 ;
        RECT  3.950 0.940 4.110 1.640 ;
        RECT  3.610 1.480 4.110 1.640 ;
        RECT  2.540 1.600 3.070 1.760 ;
        RECT  2.910 1.600 3.070 2.080 ;
        RECT  3.610 1.480 3.770 2.080 ;
        RECT  2.910 1.920 3.770 2.080 ;
        RECT  4.070 0.460 4.450 0.620 ;
        RECT  4.290 0.980 4.650 1.190 ;
        RECT  4.290 0.460 4.450 2.020 ;
        RECT  4.290 1.860 4.730 2.020 ;
        RECT  5.860 0.640 6.220 0.860 ;
        RECT  5.860 0.640 6.020 1.760 ;
        RECT  5.860 1.560 6.150 1.760 ;
        RECT  5.330 0.640 5.700 0.860 ;
        RECT  6.820 1.050 6.980 1.640 ;
        RECT  6.370 1.480 6.980 1.640 ;
        RECT  5.330 0.640 5.490 2.080 ;
        RECT  6.370 1.480 6.530 2.080 ;
        RECT  5.330 1.920 6.530 2.080 ;
        RECT  4.610 0.320 6.540 0.480 ;
        RECT  7.060 0.320 7.980 0.480 ;
        RECT  8.500 0.320 9.600 0.480 ;
        RECT  4.610 0.320 4.970 0.560 ;
        RECT  9.260 0.320 9.600 0.640 ;
        RECT  7.820 0.320 7.980 0.960 ;
        RECT  7.060 0.320 7.220 0.890 ;
        RECT  6.380 0.730 7.220 0.890 ;
        RECT  8.500 0.320 8.660 0.960 ;
        RECT  7.820 0.800 8.660 0.960 ;
        RECT  6.380 0.320 6.540 1.260 ;
        RECT  6.180 1.060 6.540 1.260 ;
        RECT  4.810 0.320 4.970 1.580 ;
        RECT  4.620 1.360 4.970 1.580 ;
        RECT  9.260 0.320 9.420 1.750 ;
        RECT  9.140 1.550 9.420 1.750 ;
        RECT  10.080 0.660 10.360 0.880 ;
        RECT  10.080 0.660 10.260 1.750 ;
        RECT  9.660 1.550 10.260 1.750 ;
        RECT  8.820 0.640 9.100 0.860 ;
        RECT  8.820 0.640 8.980 2.080 ;
        RECT  8.380 1.860 8.980 2.080 ;
        RECT  10.420 1.080 10.620 2.080 ;
        RECT  8.380 1.910 10.620 2.080 ;
        RECT  9.760 0.320 10.680 0.480 ;
        RECT  10.520 0.320 10.680 0.920 ;
        RECT  10.520 0.760 11.560 0.920 ;
        RECT  9.760 0.320 9.920 0.960 ;
        RECT  9.580 0.800 9.920 0.960 ;
        RECT  9.580 0.800 9.740 1.350 ;
        RECT  11.360 0.370 11.560 2.060 ;
        LAYER VTPH ;
        RECT  4.440 1.020 5.160 2.400 ;
        RECT  2.770 1.080 5.160 2.400 ;
        RECT  1.880 1.160 9.180 2.400 ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.880 1.180 12.000 2.400 ;
        RECT  11.310 1.140 12.000 2.400 ;
        RECT  0.000 1.230 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.020 ;
        RECT  0.000 0.000 4.440 1.080 ;
        RECT  0.000 0.000 2.770 1.140 ;
        RECT  5.160 0.000 12.000 1.140 ;
        RECT  0.400 0.000 2.770 1.160 ;
        RECT  5.160 0.000 11.310 1.160 ;
        RECT  9.180 0.000 11.310 1.180 ;
        RECT  0.400 0.000 1.880 1.230 ;
    END
END XOR4M4HM

MACRO XOR4M2HM
    CLASS CORE ;
    FOREIGN XOR4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.040 1.100 8.520 1.500 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.080 1.190 11.500 1.560 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.750 3.560 1.120 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.232  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.186  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 6.626  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.030 0.700 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.566  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 1.240 7.660 2.080 ;
        RECT  7.380 0.620 7.660 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.400 1.780 10.600 2.540 ;
        RECT  7.940 1.680 8.140 2.540 ;
        RECT  6.690 1.840 6.890 2.540 ;
        RECT  3.930 1.800 4.130 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.440 -0.140 10.640 0.600 ;
        RECT  8.140 -0.140 8.340 0.570 ;
        RECT  6.700 -0.140 6.900 0.560 ;
        RECT  3.400 -0.140 3.600 0.560 ;
        RECT  0.660 -0.140 0.860 0.750 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.650 1.620 1.760 ;
        RECT  1.420 1.540 1.700 1.760 ;
        RECT  0.140 0.470 0.340 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.860 1.280 2.060 2.080 ;
        RECT  1.100 1.920 2.060 2.080 ;
        RECT  1.820 0.640 1.980 1.120 ;
        RECT  1.820 0.960 2.380 1.120 ;
        RECT  2.220 0.960 2.380 2.080 ;
        RECT  2.220 1.920 2.750 2.080 ;
        RECT  1.020 0.320 3.060 0.480 ;
        RECT  2.900 0.320 3.060 1.440 ;
        RECT  1.020 0.320 1.180 1.350 ;
        RECT  2.900 1.280 3.450 1.440 ;
        RECT  3.290 1.280 3.450 1.780 ;
        RECT  2.140 0.640 2.740 0.800 ;
        RECT  2.540 0.640 2.740 1.760 ;
        RECT  3.950 0.940 4.110 1.640 ;
        RECT  3.610 1.480 4.110 1.640 ;
        RECT  2.540 1.600 3.070 1.760 ;
        RECT  2.910 1.600 3.070 2.100 ;
        RECT  3.610 1.480 3.770 2.100 ;
        RECT  2.910 1.940 3.770 2.100 ;
        RECT  4.070 0.460 4.450 0.620 ;
        RECT  4.290 0.980 4.650 1.190 ;
        RECT  4.290 0.460 4.450 2.020 ;
        RECT  4.290 1.860 4.730 2.020 ;
        RECT  5.860 0.620 6.220 0.840 ;
        RECT  5.860 0.620 6.020 1.760 ;
        RECT  5.860 1.560 6.150 1.760 ;
        RECT  5.330 0.620 5.700 0.840 ;
        RECT  6.800 1.060 7.000 1.640 ;
        RECT  6.370 1.480 7.000 1.640 ;
        RECT  5.330 0.620 5.490 2.080 ;
        RECT  6.370 1.480 6.530 2.080 ;
        RECT  5.330 1.920 6.530 2.080 ;
        RECT  4.610 0.300 6.540 0.460 ;
        RECT  7.060 0.300 7.980 0.460 ;
        RECT  8.500 0.300 9.660 0.460 ;
        RECT  4.610 0.300 4.970 0.560 ;
        RECT  9.260 0.300 9.660 0.560 ;
        RECT  7.820 0.300 7.980 0.890 ;
        RECT  7.060 0.300 7.220 0.880 ;
        RECT  6.380 0.720 7.220 0.880 ;
        RECT  8.500 0.300 8.660 0.890 ;
        RECT  7.820 0.730 8.660 0.890 ;
        RECT  6.380 0.300 6.540 1.260 ;
        RECT  6.240 1.060 6.540 1.260 ;
        RECT  4.810 0.300 4.970 1.580 ;
        RECT  4.620 1.360 4.970 1.580 ;
        RECT  9.260 0.300 9.420 1.750 ;
        RECT  9.140 1.550 9.420 1.750 ;
        RECT  8.820 0.620 9.100 0.840 ;
        RECT  8.820 0.620 8.980 2.080 ;
        RECT  8.380 1.860 8.980 2.080 ;
        RECT  10.040 1.100 10.240 2.080 ;
        RECT  8.380 1.910 10.240 2.080 ;
        RECT  10.960 0.370 11.160 0.920 ;
        RECT  9.580 0.760 11.160 0.920 ;
        RECT  9.580 0.760 9.740 1.420 ;
        RECT  10.760 0.760 10.920 1.940 ;
        RECT  10.760 1.740 11.200 1.940 ;
        LAYER VTPH ;
        RECT  4.440 1.020 5.180 2.400 ;
        RECT  2.770 1.080 5.180 2.400 ;
        RECT  2.770 1.140 9.180 2.400 ;
        RECT  1.880 1.160 9.180 2.400 ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.880 1.180 11.600 2.400 ;
        RECT  10.910 1.140 11.600 2.400 ;
        RECT  0.000 1.230 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.020 ;
        RECT  0.000 0.000 4.440 1.080 ;
        RECT  0.000 0.000 2.770 1.140 ;
        RECT  5.180 0.000 11.600 1.140 ;
        RECT  0.400 0.000 2.770 1.160 ;
        RECT  9.180 0.000 10.910 1.180 ;
        RECT  0.400 0.000 1.880 1.230 ;
    END
END XOR4M2HM

MACRO XOR4M1HM
    CLASS CORE ;
    FOREIGN XOR4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.080 1.190 11.500 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.040 1.100 8.520 1.500 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.850 3.750 1.120 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.180  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 7.567  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.030 0.700 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.444  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 1.240 7.660 1.870 ;
        RECT  7.380 0.620 7.660 1.870 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.400 1.780 10.600 2.540 ;
        RECT  7.940 1.680 8.140 2.540 ;
        RECT  6.690 1.720 6.890 2.540 ;
        RECT  3.930 1.800 4.130 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.440 -0.140 10.640 0.600 ;
        RECT  8.140 -0.140 8.340 0.570 ;
        RECT  6.700 -0.140 6.900 0.560 ;
        RECT  3.360 -0.140 3.640 0.630 ;
        RECT  0.660 -0.140 0.860 0.830 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.650 1.620 1.750 ;
        RECT  1.420 1.530 1.700 1.750 ;
        RECT  0.140 0.550 0.340 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.860 1.280 2.060 2.080 ;
        RECT  1.100 1.920 2.060 2.080 ;
        RECT  1.820 0.740 1.980 1.120 ;
        RECT  1.820 0.960 2.380 1.120 ;
        RECT  2.220 0.960 2.380 2.080 ;
        RECT  2.220 1.920 2.750 2.080 ;
        RECT  1.020 0.320 3.060 0.480 ;
        RECT  2.900 0.320 3.060 1.440 ;
        RECT  1.020 0.320 1.180 1.350 ;
        RECT  2.900 1.280 3.450 1.440 ;
        RECT  3.290 1.280 3.450 1.780 ;
        RECT  2.140 0.640 2.740 0.800 ;
        RECT  2.540 0.640 2.740 1.760 ;
        RECT  3.950 0.940 4.110 1.640 ;
        RECT  3.610 1.480 4.110 1.640 ;
        RECT  2.540 1.600 3.070 1.760 ;
        RECT  2.910 1.600 3.070 2.100 ;
        RECT  3.610 1.480 3.770 2.100 ;
        RECT  2.910 1.940 3.770 2.100 ;
        RECT  4.030 0.460 4.450 0.620 ;
        RECT  4.290 0.980 4.650 1.190 ;
        RECT  4.290 0.460 4.450 2.020 ;
        RECT  4.290 1.860 4.730 2.020 ;
        RECT  5.860 0.620 6.220 0.840 ;
        RECT  5.860 0.620 6.020 1.760 ;
        RECT  5.860 1.560 6.150 1.760 ;
        RECT  5.330 0.620 5.700 0.840 ;
        RECT  6.800 1.060 7.000 1.560 ;
        RECT  6.370 1.400 7.000 1.560 ;
        RECT  5.330 0.620 5.490 2.080 ;
        RECT  6.370 1.400 6.530 2.080 ;
        RECT  5.330 1.920 6.530 2.080 ;
        RECT  4.610 0.300 6.540 0.460 ;
        RECT  7.060 0.300 7.980 0.460 ;
        RECT  8.500 0.300 9.660 0.460 ;
        RECT  4.610 0.300 4.970 0.560 ;
        RECT  9.260 0.300 9.660 0.610 ;
        RECT  7.820 0.300 7.980 0.890 ;
        RECT  7.060 0.300 7.220 0.880 ;
        RECT  6.380 0.720 7.220 0.880 ;
        RECT  8.500 0.300 8.660 0.890 ;
        RECT  7.820 0.730 8.660 0.890 ;
        RECT  6.380 0.300 6.540 1.240 ;
        RECT  6.240 1.040 6.540 1.240 ;
        RECT  4.810 0.300 4.970 1.580 ;
        RECT  4.620 1.360 4.970 1.580 ;
        RECT  9.260 0.300 9.420 1.750 ;
        RECT  9.140 1.550 9.420 1.750 ;
        RECT  8.820 0.620 9.100 0.840 ;
        RECT  8.820 0.620 8.980 2.080 ;
        RECT  8.380 1.860 8.980 2.080 ;
        RECT  10.040 1.100 10.240 2.080 ;
        RECT  8.380 1.910 10.240 2.080 ;
        RECT  10.960 0.320 11.160 0.930 ;
        RECT  9.580 0.770 11.160 0.930 ;
        RECT  9.580 0.770 9.740 1.420 ;
        RECT  10.760 0.770 10.920 2.020 ;
        RECT  10.760 1.820 11.200 2.020 ;
        LAYER VTPH ;
        RECT  4.440 1.020 5.180 2.400 ;
        RECT  2.770 1.080 5.180 2.400 ;
        RECT  2.770 1.140 9.180 2.400 ;
        RECT  1.880 1.160 9.180 2.400 ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.880 1.180 11.600 2.400 ;
        RECT  10.910 1.140 11.600 2.400 ;
        RECT  0.000 1.230 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.020 ;
        RECT  0.000 0.000 4.440 1.080 ;
        RECT  0.000 0.000 2.770 1.140 ;
        RECT  5.180 0.000 11.600 1.140 ;
        RECT  0.400 0.000 2.770 1.160 ;
        RECT  9.180 0.000 10.910 1.180 ;
        RECT  0.400 0.000 1.880 1.230 ;
    END
END XOR4M1HM

MACRO XOR4M0HM
    CLASS CORE ;
    FOREIGN XOR4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.120 1.190 11.500 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.040 1.100 8.520 1.500 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.850 3.750 1.120 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.180  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 7.567  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.030 0.700 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.385  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 1.240 7.660 1.870 ;
        RECT  7.380 0.620 7.660 1.870 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.400 1.780 10.600 2.540 ;
        RECT  7.940 1.800 8.140 2.540 ;
        RECT  6.690 1.720 6.890 2.540 ;
        RECT  3.930 1.800 4.130 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.440 -0.140 10.640 0.600 ;
        RECT  8.140 -0.140 8.340 0.570 ;
        RECT  6.700 -0.140 6.900 0.560 ;
        RECT  3.440 -0.140 3.720 0.630 ;
        RECT  0.660 -0.140 0.860 0.830 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.650 1.620 1.750 ;
        RECT  1.420 1.530 1.700 1.750 ;
        RECT  0.140 0.550 0.340 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.860 1.280 2.060 2.080 ;
        RECT  1.100 1.920 2.060 2.080 ;
        RECT  1.820 0.740 1.980 1.120 ;
        RECT  1.820 0.960 2.380 1.120 ;
        RECT  2.220 0.960 2.380 2.080 ;
        RECT  2.220 1.920 2.750 2.080 ;
        RECT  1.020 0.320 3.060 0.480 ;
        RECT  2.900 0.320 3.060 1.440 ;
        RECT  1.020 0.320 1.180 1.350 ;
        RECT  2.900 1.280 3.450 1.440 ;
        RECT  3.290 1.280 3.450 1.780 ;
        RECT  2.140 0.640 2.740 0.800 ;
        RECT  2.540 0.640 2.740 1.760 ;
        RECT  3.950 0.940 4.110 1.640 ;
        RECT  3.610 1.480 4.110 1.640 ;
        RECT  2.540 1.600 3.070 1.760 ;
        RECT  2.910 1.600 3.070 2.100 ;
        RECT  3.610 1.480 3.770 2.100 ;
        RECT  2.910 1.940 3.770 2.100 ;
        RECT  4.070 0.460 4.450 0.620 ;
        RECT  4.290 0.980 4.650 1.190 ;
        RECT  4.290 0.460 4.450 2.020 ;
        RECT  4.290 1.860 4.730 2.020 ;
        RECT  5.860 0.620 6.220 0.840 ;
        RECT  5.860 0.620 6.020 1.760 ;
        RECT  5.860 1.560 6.150 1.760 ;
        RECT  5.330 0.620 5.700 0.840 ;
        RECT  6.800 1.060 7.000 1.560 ;
        RECT  6.370 1.400 7.000 1.560 ;
        RECT  5.330 0.620 5.490 2.080 ;
        RECT  6.370 1.400 6.530 2.080 ;
        RECT  5.330 1.920 6.530 2.080 ;
        RECT  4.610 0.300 6.540 0.460 ;
        RECT  7.060 0.300 7.980 0.460 ;
        RECT  8.500 0.300 9.660 0.460 ;
        RECT  4.610 0.300 4.970 0.560 ;
        RECT  9.260 0.300 9.660 0.610 ;
        RECT  7.820 0.300 7.980 0.890 ;
        RECT  7.060 0.300 7.220 0.880 ;
        RECT  6.380 0.720 7.220 0.880 ;
        RECT  8.500 0.300 8.660 0.890 ;
        RECT  7.820 0.730 8.660 0.890 ;
        RECT  6.380 0.300 6.540 1.240 ;
        RECT  6.240 1.040 6.540 1.240 ;
        RECT  4.810 0.300 4.970 1.580 ;
        RECT  4.620 1.360 4.970 1.580 ;
        RECT  9.260 0.300 9.420 1.750 ;
        RECT  9.140 1.550 9.420 1.750 ;
        RECT  8.820 0.620 9.100 0.840 ;
        RECT  8.820 0.620 8.980 2.080 ;
        RECT  8.380 1.860 8.980 2.080 ;
        RECT  10.040 1.100 10.240 2.080 ;
        RECT  8.380 1.910 10.240 2.080 ;
        RECT  11.040 0.320 11.240 0.930 ;
        RECT  9.580 0.770 11.240 0.930 ;
        RECT  9.580 0.770 9.740 1.420 ;
        RECT  10.800 0.770 10.960 2.020 ;
        RECT  10.800 1.820 11.280 2.020 ;
        LAYER VTPH ;
        RECT  4.440 1.020 5.180 2.400 ;
        RECT  2.770 1.080 5.180 2.400 ;
        RECT  2.770 1.140 9.180 2.400 ;
        RECT  1.880 1.160 9.180 2.400 ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.880 1.180 11.600 2.400 ;
        RECT  10.950 1.140 11.600 2.400 ;
        RECT  0.000 1.230 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.020 ;
        RECT  0.000 0.000 4.440 1.080 ;
        RECT  0.000 0.000 2.770 1.140 ;
        RECT  5.180 0.000 11.600 1.140 ;
        RECT  0.400 0.000 2.770 1.160 ;
        RECT  9.180 0.000 10.950 1.180 ;
        RECT  0.400 0.000 1.880 1.230 ;
    END
END XOR4M0HM

MACRO XOR3M4HM
    CLASS CORE ;
    FOREIGN XOR3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.050 3.100 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.320 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.910 1.060 6.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.513  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.900 0.480 7.100 1.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.420 1.640 7.620 2.540 ;
        RECT  6.200 1.800 6.400 2.540 ;
        RECT  4.010 1.420 4.170 2.540 ;
        RECT  2.950 2.080 3.230 2.540 ;
        RECT  0.800 1.760 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.420 -0.140 7.620 0.660 ;
        RECT  6.330 -0.140 6.530 0.560 ;
        RECT  3.990 -0.140 4.270 0.540 ;
        RECT  2.910 -0.140 3.110 0.710 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.530 0.340 0.860 ;
        RECT  0.140 0.700 0.640 0.860 ;
        RECT  1.500 1.010 1.660 1.600 ;
        RECT  0.480 1.440 1.660 1.600 ;
        RECT  0.480 0.700 0.640 1.980 ;
        RECT  0.100 1.780 0.640 1.980 ;
        RECT  1.130 0.320 2.500 0.480 ;
        RECT  2.280 0.620 2.630 0.820 ;
        RECT  1.130 0.320 1.290 1.200 ;
        RECT  0.960 1.000 1.290 1.200 ;
        RECT  2.280 0.320 2.500 1.680 ;
        RECT  2.220 1.460 2.500 1.680 ;
        RECT  1.820 0.640 2.110 0.860 ;
        RECT  1.820 0.640 1.980 2.020 ;
        RECT  2.650 1.760 3.670 1.920 ;
        RECT  1.620 1.860 2.800 2.020 ;
        RECT  3.390 1.760 3.670 2.080 ;
        RECT  3.490 0.460 3.650 1.600 ;
        RECT  3.490 0.700 4.910 0.860 ;
        RECT  4.750 0.700 4.910 1.310 ;
        RECT  3.490 0.700 3.710 1.600 ;
        RECT  3.390 1.440 3.710 1.600 ;
        RECT  5.570 0.640 5.850 0.860 ;
        RECT  4.210 1.040 4.490 1.240 ;
        RECT  4.330 1.040 4.490 2.080 ;
        RECT  5.570 0.640 5.730 2.080 ;
        RECT  4.330 1.920 5.730 2.080 ;
        RECT  5.070 0.320 6.170 0.480 ;
        RECT  6.010 0.320 6.170 0.880 ;
        RECT  6.010 0.720 6.740 0.880 ;
        RECT  6.580 0.720 6.740 1.300 ;
        RECT  5.070 0.320 5.270 1.760 ;
        RECT  4.990 1.560 5.270 1.760 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.700 2.400 ;
        RECT  3.220 1.080 4.880 2.400 ;
        RECT  6.020 1.140 8.000 2.400 ;
        RECT  0.000 1.160 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.080 ;
        RECT  0.000 0.000 3.220 1.140 ;
        RECT  4.880 0.000 8.000 1.140 ;
        RECT  1.700 0.000 3.220 1.160 ;
        RECT  4.880 0.000 6.020 1.160 ;
    END
END XOR3M4HM

MACRO XOR3M2HM
    CLASS CORE ;
    FOREIGN XOR3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.060 3.100 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.320 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.910 1.050 6.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.850 0.480 7.100 1.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.200 1.800 6.400 2.540 ;
        RECT  4.010 1.410 4.170 2.540 ;
        RECT  2.950 2.080 3.230 2.540 ;
        RECT  0.800 1.760 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.330 -0.140 6.530 0.560 ;
        RECT  3.990 -0.140 4.270 0.540 ;
        RECT  2.910 -0.140 3.110 0.620 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.550 0.340 0.860 ;
        RECT  0.140 0.700 0.640 0.860 ;
        RECT  1.500 1.010 1.660 1.600 ;
        RECT  0.480 1.440 1.660 1.600 ;
        RECT  0.480 0.700 0.640 1.980 ;
        RECT  0.100 1.780 0.640 1.980 ;
        RECT  1.130 0.300 2.500 0.460 ;
        RECT  2.280 0.600 2.630 0.800 ;
        RECT  1.130 0.300 1.290 1.200 ;
        RECT  0.960 1.000 1.290 1.200 ;
        RECT  2.280 0.300 2.500 1.680 ;
        RECT  2.220 1.460 2.500 1.680 ;
        RECT  1.820 0.620 2.110 0.840 ;
        RECT  1.820 0.620 1.980 2.020 ;
        RECT  2.650 1.760 3.670 1.920 ;
        RECT  1.620 1.860 2.800 2.020 ;
        RECT  3.390 1.760 3.670 2.080 ;
        RECT  3.490 0.460 3.650 1.600 ;
        RECT  3.490 0.700 4.910 0.860 ;
        RECT  4.750 0.700 4.910 1.310 ;
        RECT  3.490 0.700 3.710 1.600 ;
        RECT  3.390 1.440 3.710 1.600 ;
        RECT  5.570 0.620 5.850 0.840 ;
        RECT  4.210 1.040 4.490 1.240 ;
        RECT  4.330 1.040 4.490 2.080 ;
        RECT  5.570 0.620 5.730 2.080 ;
        RECT  4.330 1.920 5.730 2.080 ;
        RECT  5.070 0.300 6.170 0.460 ;
        RECT  6.010 0.300 6.170 0.880 ;
        RECT  6.010 0.720 6.690 0.880 ;
        RECT  6.530 0.720 6.690 1.300 ;
        RECT  5.070 0.300 5.270 1.760 ;
        RECT  4.990 1.560 5.270 1.760 ;
        LAYER VTPH ;
        RECT  3.250 1.080 4.880 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.080 ;
        RECT  0.000 0.000 3.250 1.140 ;
        RECT  4.880 0.000 7.200 1.140 ;
    END
END XOR3M2HM

MACRO XOR3M1HM
    CLASS CORE ;
    FOREIGN XOR3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.730 1.240 3.100 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.320 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.910 1.110 6.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.850 0.300 7.100 1.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.210 1.760 6.490 2.540 ;
        RECT  4.010 1.410 4.170 2.540 ;
        RECT  2.950 2.080 3.230 2.540 ;
        RECT  0.800 1.760 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.330 -0.140 6.530 0.580 ;
        RECT  3.990 -0.140 4.270 0.540 ;
        RECT  2.950 -0.140 3.150 0.670 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.550 0.340 0.860 ;
        RECT  0.140 0.700 0.640 0.860 ;
        RECT  1.500 1.010 1.660 1.600 ;
        RECT  0.480 1.440 1.660 1.600 ;
        RECT  0.480 0.700 0.640 1.980 ;
        RECT  0.100 1.780 0.640 1.980 ;
        RECT  1.130 0.300 2.500 0.460 ;
        RECT  2.280 0.600 2.630 0.800 ;
        RECT  1.130 0.300 1.290 1.200 ;
        RECT  0.960 1.000 1.290 1.200 ;
        RECT  2.280 0.300 2.500 1.680 ;
        RECT  2.220 1.460 2.500 1.680 ;
        RECT  1.820 0.620 2.110 0.840 ;
        RECT  1.820 0.620 1.980 2.020 ;
        RECT  2.650 1.760 3.670 1.920 ;
        RECT  1.620 1.860 2.800 2.020 ;
        RECT  3.390 1.760 3.670 2.080 ;
        RECT  3.490 0.460 3.650 1.600 ;
        RECT  3.490 0.700 4.910 0.860 ;
        RECT  4.750 0.700 4.910 1.310 ;
        RECT  3.490 0.700 3.710 1.600 ;
        RECT  3.390 1.440 3.710 1.600 ;
        RECT  5.570 0.620 5.850 0.840 ;
        RECT  4.210 1.040 4.490 1.240 ;
        RECT  4.330 1.040 4.490 2.080 ;
        RECT  5.570 0.620 5.730 2.080 ;
        RECT  4.330 1.920 5.730 2.080 ;
        RECT  5.070 0.300 6.170 0.460 ;
        RECT  6.010 0.300 6.170 0.900 ;
        RECT  6.010 0.740 6.690 0.900 ;
        RECT  6.530 0.740 6.690 1.300 ;
        RECT  5.070 0.300 5.270 1.760 ;
        RECT  4.990 1.560 5.270 1.760 ;
        LAYER VTPH ;
        RECT  3.250 1.080 4.880 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.080 ;
        RECT  0.000 0.000 3.250 1.140 ;
        RECT  4.880 0.000 7.200 1.140 ;
    END
END XOR3M1HM

MACRO XOR3M0HM
    CLASS CORE ;
    FOREIGN XOR3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.730 1.240 3.100 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.320 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.030 1.110 6.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.850 0.300 7.100 1.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.190 1.760 6.470 2.540 ;
        RECT  4.010 1.340 4.170 2.540 ;
        RECT  2.950 2.080 3.230 2.540 ;
        RECT  0.800 1.760 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.330 -0.140 6.530 0.580 ;
        RECT  3.990 -0.140 4.270 0.540 ;
        RECT  2.950 -0.140 3.150 0.670 ;
        RECT  0.740 -0.140 1.020 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.550 0.340 0.860 ;
        RECT  0.140 0.700 0.640 0.860 ;
        RECT  1.500 1.010 1.660 1.600 ;
        RECT  0.480 1.440 1.660 1.600 ;
        RECT  0.480 0.700 0.640 1.980 ;
        RECT  0.100 1.780 0.640 1.980 ;
        RECT  1.180 0.300 2.500 0.460 ;
        RECT  2.280 0.600 2.630 0.800 ;
        RECT  1.180 0.300 1.340 1.200 ;
        RECT  0.960 1.000 1.340 1.200 ;
        RECT  2.280 0.300 2.500 1.680 ;
        RECT  2.220 1.460 2.500 1.680 ;
        RECT  1.820 0.620 2.110 0.840 ;
        RECT  1.820 0.620 1.980 2.020 ;
        RECT  2.650 1.760 3.670 1.920 ;
        RECT  1.620 1.860 2.800 2.020 ;
        RECT  3.390 1.760 3.670 2.080 ;
        RECT  3.430 0.500 3.630 1.600 ;
        RECT  3.430 0.700 4.910 0.860 ;
        RECT  4.750 0.700 4.910 1.310 ;
        RECT  3.430 0.700 3.710 1.600 ;
        RECT  4.170 1.020 4.530 1.180 ;
        RECT  4.370 1.020 4.530 2.080 ;
        RECT  5.570 0.620 5.850 2.080 ;
        RECT  4.370 1.920 5.850 2.080 ;
        RECT  5.070 0.300 6.170 0.460 ;
        RECT  6.010 0.300 6.170 0.900 ;
        RECT  6.010 0.740 6.690 0.900 ;
        RECT  6.530 0.740 6.690 1.300 ;
        RECT  5.070 0.300 5.270 1.760 ;
        RECT  4.990 1.560 5.270 1.760 ;
        LAYER VTPH ;
        RECT  3.250 1.080 4.880 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.080 ;
        RECT  0.000 0.000 3.250 1.140 ;
        RECT  4.880 0.000 7.200 1.140 ;
    END
END XOR3M0HM

MACRO XOR2M8HM
    CLASS CORE ;
    FOREIGN XOR2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 0.840 4.400 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 1.120 1.220 ;
        RECT  0.100 0.840 0.300 1.220 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 0.420 6.300 2.100 ;
        RECT  5.080 1.440 6.300 1.640 ;
        RECT  5.080 0.660 6.300 0.860 ;
        RECT  5.080 1.440 5.280 2.100 ;
        RECT  5.080 0.420 5.280 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.640 1.720 6.840 2.540 ;
        RECT  5.600 1.800 5.800 2.540 ;
        RECT  4.580 1.800 4.780 2.540 ;
        RECT  1.160 1.770 1.360 2.540 ;
        RECT  0.140 1.720 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.640 -0.140 6.840 0.680 ;
        RECT  5.560 -0.140 5.840 0.500 ;
        RECT  4.560 -0.140 4.760 0.680 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.720 0.380 1.880 1.160 ;
        RECT  1.840 1.000 2.000 1.780 ;
        RECT  0.680 0.380 0.840 0.820 ;
        RECT  0.680 0.660 1.540 0.820 ;
        RECT  2.780 0.620 3.080 0.840 ;
        RECT  1.380 0.660 1.540 1.610 ;
        RECT  0.660 1.450 1.680 1.610 ;
        RECT  1.520 1.450 1.680 2.100 ;
        RECT  0.660 1.450 0.860 2.100 ;
        RECT  2.920 0.620 3.080 2.100 ;
        RECT  1.520 1.940 3.080 2.100 ;
        RECT  3.760 0.500 4.320 0.660 ;
        RECT  3.760 0.500 3.920 1.780 ;
        RECT  3.760 1.500 4.100 1.780 ;
        RECT  2.360 0.300 3.600 0.460 ;
        RECT  2.140 0.500 2.520 0.660 ;
        RECT  4.760 1.060 5.900 1.220 ;
        RECT  4.760 1.060 4.920 1.640 ;
        RECT  4.260 1.480 4.920 1.640 ;
        RECT  2.360 0.300 2.520 1.780 ;
        RECT  3.440 0.300 3.600 2.100 ;
        RECT  4.260 1.480 4.420 2.100 ;
        RECT  3.440 1.940 4.420 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END XOR2M8HM

MACRO XOR2M6HM
    CLASS CORE ;
    FOREIGN XOR2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.650 0.840 3.940 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.120 1.240 ;
        RECT  0.100 0.840 0.300 1.240 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.680 1.440 5.900 2.100 ;
        RECT  5.700 0.420 5.900 2.100 ;
        RECT  4.620 0.660 5.900 0.860 ;
        RECT  5.680 0.420 5.900 0.860 ;
        RECT  4.620 1.440 5.900 1.640 ;
        RECT  4.620 1.440 4.820 2.100 ;
        RECT  4.620 0.420 4.820 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.140 1.800 5.340 2.540 ;
        RECT  4.120 1.780 4.320 2.540 ;
        RECT  1.160 1.770 1.360 2.540 ;
        RECT  0.140 1.720 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.380 0.500 ;
        RECT  4.100 -0.140 4.300 0.680 ;
        RECT  1.160 -0.140 1.360 0.600 ;
        RECT  0.140 -0.140 0.340 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.840 0.620 2.060 0.900 ;
        RECT  1.840 0.620 2.000 1.930 ;
        RECT  1.620 1.770 2.000 1.930 ;
        RECT  1.520 0.300 3.140 0.460 ;
        RECT  0.680 0.340 0.840 0.920 ;
        RECT  1.520 0.300 1.680 0.920 ;
        RECT  0.680 0.760 1.680 0.920 ;
        RECT  1.380 0.760 1.540 1.610 ;
        RECT  0.660 1.450 1.540 1.610 ;
        RECT  2.980 0.300 3.140 1.780 ;
        RECT  2.700 1.620 3.140 1.780 ;
        RECT  0.660 1.450 0.860 1.940 ;
        RECT  3.300 0.500 3.860 0.660 ;
        RECT  3.300 0.500 3.460 1.780 ;
        RECT  3.300 1.500 3.640 1.780 ;
        RECT  2.240 0.660 2.720 0.820 ;
        RECT  4.140 1.060 5.440 1.220 ;
        RECT  4.140 1.060 4.300 1.620 ;
        RECT  3.800 1.460 4.300 1.620 ;
        RECT  2.240 0.660 2.400 2.100 ;
        RECT  3.800 1.460 3.960 2.100 ;
        RECT  2.240 1.940 3.960 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.480 2.400 ;
        RECT  3.500 1.140 6.000 2.400 ;
        RECT  0.000 1.200 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
        RECT  1.480 0.000 3.500 1.200 ;
    END
END XOR2M6HM

MACRO XOR2M4HM
    CLASS CORE ;
    FOREIGN XOR2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 0.840 3.100 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.620 1.360 4.300 1.560 ;
        RECT  4.100 0.660 4.300 1.560 ;
        RECT  3.620 0.660 4.300 0.860 ;
        RECT  3.620 1.360 3.820 2.100 ;
        RECT  3.620 0.420 3.820 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.140 1.720 4.340 2.540 ;
        RECT  3.120 1.760 3.320 2.540 ;
        RECT  0.640 1.770 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.100 -0.140 4.380 0.500 ;
        RECT  3.100 -0.140 3.300 0.680 ;
        RECT  0.640 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.600 0.840 ;
        RECT  1.320 0.620 1.480 1.780 ;
        RECT  0.100 0.450 0.380 0.650 ;
        RECT  0.100 0.450 0.260 1.990 ;
        RECT  0.100 1.440 1.160 1.600 ;
        RECT  1.000 1.440 1.160 2.100 ;
        RECT  0.100 1.440 0.320 1.990 ;
        RECT  1.640 1.000 1.800 2.100 ;
        RECT  1.000 1.940 1.800 2.100 ;
        RECT  1.000 0.300 2.520 0.460 ;
        RECT  2.360 0.520 2.860 0.680 ;
        RECT  1.000 0.300 1.160 1.280 ;
        RECT  0.900 1.000 1.160 1.280 ;
        RECT  2.360 0.300 2.520 1.780 ;
        RECT  2.360 1.500 2.640 1.780 ;
        RECT  1.920 0.620 2.200 0.840 ;
        RECT  3.300 1.040 3.900 1.200 ;
        RECT  3.300 1.040 3.460 1.600 ;
        RECT  2.800 1.440 3.460 1.600 ;
        RECT  1.960 0.620 2.120 2.100 ;
        RECT  2.800 1.440 2.960 2.100 ;
        RECT  1.960 1.940 2.960 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END XOR2M4HM

MACRO XOR2M3HM
    CLASS CORE ;
    FOREIGN XOR2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 0.840 3.100 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.620 1.360 4.300 1.560 ;
        RECT  4.100 0.660 4.300 1.560 ;
        RECT  3.620 0.660 4.300 0.860 ;
        RECT  3.620 1.360 3.820 1.980 ;
        RECT  3.620 0.340 3.820 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.140 1.720 4.340 2.540 ;
        RECT  3.120 1.760 3.320 2.540 ;
        RECT  0.640 1.770 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.100 -0.140 4.380 0.500 ;
        RECT  3.100 -0.140 3.300 0.680 ;
        RECT  0.640 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.600 0.840 ;
        RECT  1.320 0.620 1.480 1.780 ;
        RECT  0.100 0.450 0.380 0.650 ;
        RECT  0.100 0.450 0.260 1.990 ;
        RECT  0.100 1.440 1.160 1.600 ;
        RECT  1.000 1.440 1.160 2.100 ;
        RECT  0.100 1.440 0.320 1.990 ;
        RECT  1.640 1.000 1.800 2.100 ;
        RECT  1.000 1.940 1.800 2.100 ;
        RECT  1.000 0.300 2.520 0.460 ;
        RECT  2.360 0.520 2.860 0.680 ;
        RECT  1.000 0.300 1.160 1.280 ;
        RECT  0.900 1.000 1.160 1.280 ;
        RECT  2.360 0.300 2.520 1.780 ;
        RECT  2.360 1.500 2.640 1.780 ;
        RECT  1.920 0.620 2.200 0.840 ;
        RECT  3.300 1.040 3.900 1.200 ;
        RECT  3.300 1.040 3.460 1.600 ;
        RECT  2.800 1.440 3.460 1.600 ;
        RECT  1.960 0.620 2.120 2.100 ;
        RECT  2.800 1.440 2.960 2.100 ;
        RECT  1.960 1.940 2.960 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END XOR2M3HM

MACRO XOR2M2HM
    CLASS CORE ;
    FOREIGN XOR2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.640 0.420 3.900 2.100 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 0.840 3.100 1.280 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.120 1.760 3.320 2.540 ;
        RECT  0.640 1.770 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.100 -0.140 3.300 0.680 ;
        RECT  0.640 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.600 0.840 ;
        RECT  1.320 0.620 1.480 1.780 ;
        RECT  0.100 0.450 0.380 0.650 ;
        RECT  0.100 0.450 0.260 1.990 ;
        RECT  0.100 1.440 1.160 1.600 ;
        RECT  1.000 1.440 1.160 2.100 ;
        RECT  0.100 1.440 0.320 1.990 ;
        RECT  1.640 1.000 1.800 2.100 ;
        RECT  1.000 1.940 1.800 2.100 ;
        RECT  1.000 0.300 2.520 0.460 ;
        RECT  2.360 0.520 2.860 0.680 ;
        RECT  1.000 0.300 1.160 1.280 ;
        RECT  0.900 1.000 1.160 1.280 ;
        RECT  2.360 0.300 2.520 1.780 ;
        RECT  2.360 1.500 2.640 1.780 ;
        RECT  1.920 0.620 2.200 0.840 ;
        RECT  3.300 0.960 3.460 1.600 ;
        RECT  2.800 1.440 3.460 1.600 ;
        RECT  1.960 0.620 2.120 2.100 ;
        RECT  2.800 1.440 2.960 2.100 ;
        RECT  1.960 1.940 2.960 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END XOR2M2HM

MACRO XOR2M1HM
    CLASS CORE ;
    FOREIGN XOR2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.640 0.420 3.900 1.940 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 0.840 3.100 1.280 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.120 1.760 3.320 2.540 ;
        RECT  0.640 1.770 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.100 -0.140 3.300 0.680 ;
        RECT  0.640 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.600 0.840 ;
        RECT  1.320 0.620 1.480 1.780 ;
        RECT  0.100 0.450 0.380 0.650 ;
        RECT  0.100 0.450 0.260 1.990 ;
        RECT  0.100 1.440 1.160 1.600 ;
        RECT  1.000 1.440 1.160 2.100 ;
        RECT  0.100 1.440 0.320 1.990 ;
        RECT  1.640 1.000 1.800 2.100 ;
        RECT  1.000 1.940 1.800 2.100 ;
        RECT  1.000 0.300 2.520 0.460 ;
        RECT  2.360 0.520 2.860 0.680 ;
        RECT  1.000 0.300 1.160 1.280 ;
        RECT  0.900 1.000 1.160 1.280 ;
        RECT  2.360 0.300 2.520 1.780 ;
        RECT  2.360 1.500 2.640 1.780 ;
        RECT  1.920 0.620 2.200 0.840 ;
        RECT  3.300 0.960 3.460 1.600 ;
        RECT  2.800 1.440 3.460 1.600 ;
        RECT  1.960 0.620 2.120 2.100 ;
        RECT  2.800 1.440 2.960 2.100 ;
        RECT  1.960 1.940 2.960 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END XOR2M1HM

MACRO XOR2M0HM
    CLASS CORE ;
    FOREIGN XOR2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.640 0.400 3.900 1.940 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 0.840 3.100 1.280 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.120 1.760 3.320 2.540 ;
        RECT  0.640 1.770 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.100 -0.140 3.300 0.680 ;
        RECT  0.640 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.600 0.840 ;
        RECT  1.320 0.620 1.480 1.780 ;
        RECT  0.100 0.450 0.380 0.650 ;
        RECT  0.100 0.450 0.260 1.990 ;
        RECT  0.100 1.440 1.160 1.600 ;
        RECT  1.000 1.440 1.160 2.100 ;
        RECT  0.100 1.440 0.320 1.990 ;
        RECT  1.640 1.000 1.800 2.100 ;
        RECT  1.000 1.940 1.800 2.100 ;
        RECT  1.000 0.300 2.520 0.460 ;
        RECT  2.360 0.460 2.860 0.620 ;
        RECT  1.000 0.300 1.160 1.280 ;
        RECT  0.900 1.000 1.160 1.280 ;
        RECT  2.360 0.300 2.520 1.780 ;
        RECT  2.360 1.500 2.640 1.780 ;
        RECT  1.920 0.620 2.200 0.840 ;
        RECT  3.300 0.960 3.460 1.600 ;
        RECT  2.800 1.440 3.460 1.600 ;
        RECT  1.960 0.620 2.120 2.100 ;
        RECT  2.800 1.440 2.960 2.100 ;
        RECT  1.960 1.940 2.960 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END XOR2M0HM

MACRO XNR4M4HM
    CLASS CORE ;
    FOREIGN XNR4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER ME1  ;
        ANTENNAGATEAREA 0.132  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.348  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.980 1.240 8.180 1.440 ;
        LAYER ME2 ;
        RECT  7.880 1.240 8.300 1.560 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  7.970 1.070 8.190 1.700 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.484  LAYER ME1  ;
        ANTENNADIFFAREA 0.484  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.270 1.240 7.470 1.440 ;
        LAYER ME2 ;
        RECT  7.270 0.840 7.510 1.560 ;
        LAYER ME1 ;
        RECT  7.080 1.140 7.470 1.600 ;
        RECT  7.080 0.440 7.240 1.600 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.460 1.140 10.750 1.610 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.900 3.320 1.280 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.320 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.210 1.760 10.370 2.540 ;
        RECT  7.650 2.080 7.960 2.540 ;
        RECT  6.530 2.080 6.810 2.540 ;
        RECT  4.240 1.760 4.400 2.540 ;
        RECT  3.260 2.080 3.550 2.540 ;
        RECT  0.590 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.260 -0.140 10.540 0.560 ;
        RECT  7.560 -0.140 7.760 0.590 ;
        RECT  6.520 -0.140 6.680 0.420 ;
        RECT  4.200 -0.140 4.360 0.820 ;
        RECT  3.060 -0.140 3.330 0.660 ;
        RECT  0.590 -0.140 0.840 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.650 1.600 0.810 ;
        RECT  1.320 0.650 1.540 1.760 ;
        RECT  0.080 0.420 0.390 0.660 ;
        RECT  0.080 0.420 0.240 2.050 ;
        RECT  0.080 1.480 1.160 1.640 ;
        RECT  1.000 1.480 1.160 2.100 ;
        RECT  0.080 1.480 0.320 2.050 ;
        RECT  1.760 1.050 1.920 2.100 ;
        RECT  1.000 1.940 1.920 2.100 ;
        RECT  1.000 0.330 2.810 0.490 ;
        RECT  2.520 0.330 2.810 0.740 ;
        RECT  1.000 0.330 1.160 1.310 ;
        RECT  0.870 1.030 1.160 1.310 ;
        RECT  2.520 0.330 2.680 1.600 ;
        RECT  2.520 1.440 3.030 1.600 ;
        RECT  1.920 0.650 2.280 0.810 ;
        RECT  2.940 1.760 4.030 1.920 ;
        RECT  2.080 0.650 2.280 2.100 ;
        RECT  2.940 1.760 3.100 2.100 ;
        RECT  2.080 1.940 3.100 2.100 ;
        RECT  3.740 1.760 4.030 2.100 ;
        RECT  4.840 0.650 5.130 0.870 ;
        RECT  4.880 0.650 5.130 1.780 ;
        RECT  5.290 1.050 5.720 1.330 ;
        RECT  3.520 0.450 3.810 1.600 ;
        RECT  3.520 1.440 4.720 1.600 ;
        RECT  4.560 1.440 4.720 2.100 ;
        RECT  5.290 1.050 5.450 2.100 ;
        RECT  4.560 1.940 5.450 2.100 ;
        RECT  5.330 0.670 6.040 0.830 ;
        RECT  5.880 0.940 6.580 1.220 ;
        RECT  5.880 0.670 6.040 1.790 ;
        RECT  5.680 1.490 6.040 1.790 ;
        RECT  7.920 0.300 9.000 0.460 ;
        RECT  4.520 0.330 6.360 0.490 ;
        RECT  6.200 0.330 6.360 0.740 ;
        RECT  6.200 0.580 6.900 0.740 ;
        RECT  7.920 0.300 8.100 0.910 ;
        RECT  7.650 0.750 8.100 0.910 ;
        RECT  4.520 0.330 4.680 1.280 ;
        RECT  4.360 1.070 4.720 1.280 ;
        RECT  8.800 0.300 9.000 1.750 ;
        RECT  6.740 0.580 6.900 1.920 ;
        RECT  6.270 1.450 6.900 1.920 ;
        RECT  7.650 0.750 7.810 1.920 ;
        RECT  6.270 1.760 7.810 1.920 ;
        RECT  9.480 0.620 9.770 0.940 ;
        RECT  9.480 0.620 9.730 1.730 ;
        RECT  9.320 1.570 9.730 1.730 ;
        RECT  8.260 0.620 8.540 0.920 ;
        RECT  9.890 1.090 10.090 1.440 ;
        RECT  8.360 0.620 8.540 2.070 ;
        RECT  8.170 1.860 8.540 2.070 ;
        RECT  9.890 1.090 10.050 2.070 ;
        RECT  8.170 1.910 10.050 2.070 ;
        RECT  9.160 0.300 10.100 0.460 ;
        RECT  9.940 0.300 10.100 0.920 ;
        RECT  10.770 0.520 11.080 0.920 ;
        RECT  9.940 0.760 11.080 0.920 ;
        RECT  9.160 0.300 9.320 1.360 ;
        RECT  10.920 0.520 11.080 2.060 ;
        RECT  10.610 1.830 11.080 2.060 ;
        LAYER VTPH ;
        RECT  6.450 1.080 8.030 2.400 ;
        RECT  0.000 1.140 1.050 2.400 ;
        RECT  2.470 1.080 4.080 2.400 ;
        RECT  0.000 1.170 4.080 2.400 ;
        RECT  6.450 1.150 9.210 2.400 ;
        RECT  10.400 1.140 11.200 2.400 ;
        RECT  0.000 1.190 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.080 ;
        RECT  0.000 0.000 2.470 1.140 ;
        RECT  8.030 0.000 11.200 1.140 ;
        RECT  8.030 0.000 10.400 1.150 ;
        RECT  1.050 0.000 2.470 1.170 ;
        RECT  4.080 0.000 6.450 1.190 ;
        RECT  9.210 0.000 10.400 1.190 ;
    END
END XNR4M4HM

MACRO XNR4M2HM
    CLASS CORE ;
    FOREIGN XNR4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.394  LAYER ME1  ;
        ANTENNADIFFAREA 0.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.870 1.240 7.070 1.440 ;
        LAYER ME2 ;
        RECT  6.870 0.840 7.110 1.560 ;
        LAYER ME1 ;
        RECT  6.750 1.140 7.070 1.600 ;
        RECT  6.750 0.440 6.910 1.600 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER ME1  ;
        ANTENNAGATEAREA 0.132  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.348  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.650 1.240 7.850 1.440 ;
        LAYER ME2 ;
        RECT  7.650 0.840 7.970 1.560 ;
        LAYER ME1 ;
        RECT  7.640 1.070 7.860 1.700 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.060 1.140 10.350 1.610 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.900 3.320 1.280 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.320 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  9.810 1.760 9.970 2.540 ;
        RECT  7.320 2.080 7.630 2.540 ;
        RECT  4.240 1.760 4.400 2.540 ;
        RECT  3.260 2.080 3.550 2.540 ;
        RECT  0.590 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  9.660 -0.140 9.940 0.560 ;
        RECT  7.230 -0.140 7.430 0.590 ;
        RECT  4.200 -0.140 4.360 0.820 ;
        RECT  3.060 -0.140 3.330 0.660 ;
        RECT  0.590 -0.140 0.840 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.650 1.600 0.810 ;
        RECT  1.320 0.650 1.540 1.760 ;
        RECT  0.080 0.420 0.390 0.660 ;
        RECT  0.080 0.420 0.240 2.050 ;
        RECT  0.080 1.480 1.160 1.640 ;
        RECT  1.000 1.480 1.160 2.100 ;
        RECT  0.080 1.480 0.320 2.050 ;
        RECT  1.760 1.050 1.920 2.100 ;
        RECT  1.000 1.940 1.920 2.100 ;
        RECT  1.000 0.330 2.810 0.490 ;
        RECT  2.520 0.330 2.810 0.740 ;
        RECT  1.000 0.330 1.160 1.310 ;
        RECT  0.870 1.030 1.160 1.310 ;
        RECT  2.520 0.330 2.680 1.600 ;
        RECT  2.520 1.440 3.030 1.600 ;
        RECT  1.920 0.650 2.280 0.810 ;
        RECT  2.940 1.760 4.030 1.920 ;
        RECT  2.080 0.650 2.280 2.100 ;
        RECT  2.940 1.760 3.100 2.100 ;
        RECT  2.080 1.940 3.100 2.100 ;
        RECT  3.740 1.760 4.030 2.100 ;
        RECT  4.840 0.650 5.130 0.870 ;
        RECT  4.880 0.650 5.130 1.780 ;
        RECT  5.290 1.050 5.720 1.330 ;
        RECT  3.520 0.450 3.810 1.600 ;
        RECT  3.520 1.440 4.720 1.600 ;
        RECT  4.560 1.440 4.720 2.100 ;
        RECT  5.290 1.050 5.450 2.100 ;
        RECT  4.560 1.940 5.450 2.100 ;
        RECT  5.330 0.670 6.040 0.830 ;
        RECT  5.880 1.000 6.250 1.280 ;
        RECT  5.880 0.670 6.040 2.080 ;
        RECT  5.720 1.730 6.040 2.080 ;
        RECT  7.590 0.300 8.670 0.460 ;
        RECT  4.520 0.330 6.570 0.490 ;
        RECT  7.590 0.300 7.770 0.910 ;
        RECT  7.320 0.750 7.770 0.910 ;
        RECT  4.520 0.330 4.680 1.280 ;
        RECT  4.360 1.020 4.680 1.280 ;
        RECT  8.470 0.300 8.670 1.750 ;
        RECT  6.410 0.330 6.570 1.920 ;
        RECT  6.410 1.760 7.480 1.920 ;
        RECT  7.320 0.750 7.480 1.920 ;
        RECT  6.210 1.770 6.520 2.080 ;
        RECT  7.930 0.620 8.210 0.920 ;
        RECT  9.490 1.090 9.690 1.440 ;
        RECT  8.030 0.620 8.210 2.070 ;
        RECT  7.840 1.860 8.210 2.070 ;
        RECT  9.490 1.090 9.650 2.070 ;
        RECT  7.840 1.910 9.650 2.070 ;
        RECT  10.370 0.520 10.680 0.920 ;
        RECT  8.830 0.760 10.680 0.920 ;
        RECT  8.830 0.760 8.990 1.360 ;
        RECT  10.520 0.520 10.680 2.060 ;
        RECT  10.210 1.830 10.680 2.060 ;
        LAYER VTPH ;
        RECT  6.450 1.080 7.700 2.400 ;
        RECT  0.000 1.140 1.050 2.400 ;
        RECT  2.470 1.080 4.080 2.400 ;
        RECT  0.000 1.170 4.080 2.400 ;
        RECT  6.450 1.150 8.880 2.400 ;
        RECT  10.000 1.140 10.800 2.400 ;
        RECT  0.000 1.190 10.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.800 1.080 ;
        RECT  0.000 0.000 2.470 1.140 ;
        RECT  7.700 0.000 10.800 1.140 ;
        RECT  7.700 0.000 10.000 1.150 ;
        RECT  1.050 0.000 2.470 1.170 ;
        RECT  4.080 0.000 6.450 1.190 ;
        RECT  8.880 0.000 10.000 1.190 ;
    END
END XNR4M2HM

MACRO XNR4M1HM
    CLASS CORE ;
    FOREIGN XNR4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        ANTENNADIFFAREA 0.296  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.240 7.100 1.440 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.140 1.560 ;
        LAYER ME1 ;
        RECT  6.820 1.140 7.140 1.600 ;
        RECT  6.820 0.370 6.980 1.600 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.385  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.730 1.240 7.930 1.440 ;
        LAYER ME2 ;
        RECT  7.700 0.840 7.930 1.560 ;
        LAYER ME1 ;
        RECT  7.710 1.070 7.930 1.700 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.155  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.040 1.140 10.350 1.610 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.900 3.390 1.280 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.320 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  9.810 1.760 9.970 2.540 ;
        RECT  7.390 2.080 7.700 2.540 ;
        RECT  4.310 1.760 4.470 2.540 ;
        RECT  3.260 2.080 3.620 2.540 ;
        RECT  0.590 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  9.660 -0.140 9.940 0.560 ;
        RECT  7.300 -0.140 7.500 0.590 ;
        RECT  4.270 -0.140 4.430 0.820 ;
        RECT  3.130 -0.140 3.330 0.680 ;
        RECT  0.590 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.650 1.600 0.810 ;
        RECT  1.320 0.650 1.540 1.760 ;
        RECT  0.080 0.420 0.390 0.660 ;
        RECT  0.080 0.420 0.240 2.050 ;
        RECT  0.080 1.480 1.160 1.640 ;
        RECT  1.000 1.480 1.160 2.100 ;
        RECT  0.080 1.480 0.320 2.050 ;
        RECT  1.760 1.050 1.920 2.100 ;
        RECT  1.000 1.940 1.920 2.100 ;
        RECT  1.000 0.330 2.810 0.490 ;
        RECT  2.520 0.330 2.810 0.740 ;
        RECT  1.000 0.330 1.160 1.310 ;
        RECT  0.870 1.030 1.160 1.310 ;
        RECT  2.520 0.330 2.680 1.600 ;
        RECT  2.520 1.440 3.030 1.600 ;
        RECT  1.920 0.650 2.280 0.810 ;
        RECT  2.940 1.760 4.100 1.920 ;
        RECT  2.080 0.650 2.280 2.100 ;
        RECT  2.940 1.760 3.100 2.100 ;
        RECT  2.080 1.940 3.100 2.100 ;
        RECT  3.810 1.760 4.100 2.100 ;
        RECT  4.910 0.650 5.200 0.870 ;
        RECT  4.950 0.650 5.200 1.780 ;
        RECT  5.360 1.050 5.790 1.330 ;
        RECT  3.590 0.450 3.880 1.600 ;
        RECT  3.590 1.440 4.790 1.600 ;
        RECT  4.630 1.440 4.790 2.100 ;
        RECT  5.360 1.050 5.520 2.100 ;
        RECT  4.630 1.940 5.520 2.100 ;
        RECT  5.400 0.670 6.110 0.830 ;
        RECT  5.950 1.000 6.320 1.280 ;
        RECT  5.950 0.670 6.110 2.080 ;
        RECT  5.790 1.730 6.110 2.080 ;
        RECT  7.660 0.300 8.740 0.460 ;
        RECT  4.590 0.330 6.640 0.490 ;
        RECT  7.660 0.300 7.840 0.910 ;
        RECT  7.390 0.750 7.840 0.910 ;
        RECT  4.590 0.330 4.750 1.280 ;
        RECT  4.430 1.020 4.750 1.280 ;
        RECT  8.540 0.300 8.740 1.750 ;
        RECT  6.480 0.330 6.640 1.920 ;
        RECT  6.480 1.760 7.550 1.920 ;
        RECT  7.390 0.750 7.550 1.920 ;
        RECT  6.280 1.770 6.590 2.080 ;
        RECT  8.000 0.620 8.280 0.920 ;
        RECT  8.100 0.620 8.280 2.070 ;
        RECT  7.910 1.860 8.280 2.070 ;
        RECT  9.400 1.040 9.650 2.070 ;
        RECT  7.910 1.910 9.650 2.070 ;
        RECT  10.370 0.520 10.700 0.880 ;
        RECT  8.900 0.720 10.700 0.880 ;
        RECT  8.900 0.720 9.060 1.360 ;
        RECT  10.520 0.520 10.700 2.060 ;
        RECT  10.210 1.830 10.700 2.060 ;
        LAYER VTPH ;
        RECT  6.520 1.080 7.770 2.400 ;
        RECT  0.000 1.140 1.050 2.400 ;
        RECT  2.460 1.080 4.150 2.400 ;
        RECT  0.000 1.170 4.150 2.400 ;
        RECT  6.520 1.150 8.950 2.400 ;
        RECT  10.000 1.140 10.800 2.400 ;
        RECT  0.000 1.190 10.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.800 1.080 ;
        RECT  0.000 0.000 2.460 1.140 ;
        RECT  7.770 0.000 10.800 1.140 ;
        RECT  7.770 0.000 10.000 1.150 ;
        RECT  1.050 0.000 2.460 1.170 ;
        RECT  4.150 0.000 6.520 1.190 ;
        RECT  8.950 0.000 10.000 1.190 ;
    END
END XNR4M1HM

MACRO XNR4M0HM
    CLASS CORE ;
    FOREIGN XNR4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        ANTENNADIFFAREA 0.235  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.240 7.100 1.440 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.140 1.560 ;
        LAYER ME1 ;
        RECT  6.820 0.300 7.140 1.600 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        ANTENNAGATEAREA 0.060  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.367  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.730 1.240 7.930 1.440 ;
        LAYER ME2 ;
        RECT  7.700 0.840 7.930 1.560 ;
        LAYER ME1 ;
        RECT  7.710 1.070 7.930 1.700 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.040 1.140 10.350 1.610 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.061  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.900 3.390 1.280 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.320 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  9.810 1.760 9.970 2.540 ;
        RECT  7.390 2.080 7.700 2.540 ;
        RECT  4.310 1.760 4.470 2.540 ;
        RECT  3.260 2.080 3.620 2.540 ;
        RECT  0.590 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  9.610 -0.140 9.890 0.560 ;
        RECT  7.300 -0.140 7.500 0.590 ;
        RECT  4.270 -0.140 4.430 0.820 ;
        RECT  3.130 -0.140 3.340 0.680 ;
        RECT  0.590 -0.140 0.840 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.650 1.600 0.810 ;
        RECT  1.320 0.650 1.540 1.760 ;
        RECT  0.080 0.420 0.390 0.660 ;
        RECT  0.080 0.420 0.240 2.050 ;
        RECT  0.080 1.480 1.160 1.640 ;
        RECT  1.000 1.480 1.160 2.100 ;
        RECT  0.080 1.480 0.320 2.050 ;
        RECT  1.760 1.050 1.920 2.100 ;
        RECT  1.000 1.940 1.920 2.100 ;
        RECT  1.000 0.330 2.810 0.490 ;
        RECT  2.520 0.330 2.810 0.740 ;
        RECT  1.000 0.330 1.160 1.310 ;
        RECT  0.870 1.030 1.160 1.310 ;
        RECT  2.520 0.330 2.680 1.600 ;
        RECT  2.520 1.440 3.030 1.600 ;
        RECT  1.920 0.650 2.280 0.810 ;
        RECT  2.940 1.760 4.110 1.920 ;
        RECT  2.080 0.650 2.280 2.100 ;
        RECT  2.940 1.760 3.100 2.100 ;
        RECT  2.080 1.940 3.100 2.100 ;
        RECT  3.820 1.760 4.110 2.100 ;
        RECT  4.910 0.650 5.200 0.870 ;
        RECT  4.950 0.650 5.200 1.780 ;
        RECT  5.360 1.050 5.790 1.330 ;
        RECT  3.570 0.450 3.860 1.600 ;
        RECT  3.570 1.440 4.790 1.600 ;
        RECT  4.630 1.440 4.790 2.100 ;
        RECT  5.360 1.050 5.520 2.100 ;
        RECT  4.630 1.940 5.520 2.100 ;
        RECT  5.400 0.670 6.110 0.830 ;
        RECT  5.950 1.000 6.320 1.280 ;
        RECT  5.950 0.670 6.110 2.080 ;
        RECT  5.790 1.730 6.110 2.080 ;
        RECT  7.660 0.300 8.740 0.460 ;
        RECT  4.590 0.330 6.640 0.490 ;
        RECT  7.660 0.300 7.840 0.910 ;
        RECT  7.390 0.750 7.840 0.910 ;
        RECT  4.590 0.330 4.750 1.280 ;
        RECT  4.430 1.020 4.750 1.280 ;
        RECT  8.540 0.300 8.740 1.750 ;
        RECT  6.480 0.330 6.640 1.920 ;
        RECT  6.480 1.760 7.550 1.920 ;
        RECT  7.390 0.750 7.550 1.920 ;
        RECT  6.280 1.770 6.590 2.080 ;
        RECT  8.000 0.620 8.280 0.920 ;
        RECT  8.100 0.620 8.280 2.070 ;
        RECT  7.910 1.860 8.280 2.070 ;
        RECT  9.400 1.040 9.650 2.070 ;
        RECT  7.910 1.910 9.650 2.070 ;
        RECT  10.370 0.520 10.700 0.880 ;
        RECT  8.900 0.720 10.700 0.880 ;
        RECT  8.900 0.720 9.060 1.360 ;
        RECT  10.520 0.520 10.700 2.060 ;
        RECT  10.210 1.830 10.700 2.060 ;
        LAYER VTPH ;
        RECT  6.520 1.080 7.770 2.400 ;
        RECT  0.000 1.140 1.050 2.400 ;
        RECT  2.460 1.080 4.150 2.400 ;
        RECT  0.000 1.170 4.150 2.400 ;
        RECT  6.520 1.150 8.950 2.400 ;
        RECT  10.000 1.140 10.800 2.400 ;
        RECT  0.000 1.190 10.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.800 1.080 ;
        RECT  0.000 0.000 2.460 1.140 ;
        RECT  7.770 0.000 10.800 1.140 ;
        RECT  7.770 0.000 10.000 1.150 ;
        RECT  1.050 0.000 2.460 1.170 ;
        RECT  4.150 0.000 6.520 1.190 ;
        RECT  8.950 0.000 10.000 1.190 ;
    END
END XNR4M0HM

MACRO XNR3M4HM
    CLASS CORE ;
    FOREIGN XNR3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        ANTENNAGATEAREA 0.146  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.481  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 0.680 3.100 0.880 ;
        LAYER ME2 ;
        RECT  2.900 0.440 3.100 1.160 ;
        LAYER ME1 ;
        RECT  2.490 0.620 3.140 0.950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.446  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.940 1.240 8.300 1.560 ;
        RECT  7.940 0.480 8.170 1.560 ;
        RECT  7.940 0.480 8.160 2.100 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.204  LAYER ME1  ;
        ANTENNAGATEAREA 0.204  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.810  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.310 1.440 6.510 1.640 ;
        LAYER ME2 ;
        RECT  6.100 1.380 6.510 1.960 ;
        LAYER ME1 ;
        RECT  6.260 1.380 6.570 1.780 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.460 1.470 8.660 2.540 ;
        RECT  7.440 1.430 7.600 2.540 ;
        RECT  3.940 1.440 4.100 2.540 ;
        RECT  0.660 1.800 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.460 -0.140 8.660 0.760 ;
        RECT  7.440 -0.140 7.600 0.800 ;
        RECT  3.880 -0.140 4.080 0.620 ;
        RECT  0.660 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.620 1.620 1.700 ;
        RECT  1.020 0.300 2.900 0.460 ;
        RECT  0.140 1.480 1.180 1.640 ;
        RECT  1.020 0.300 1.180 2.020 ;
        RECT  1.020 1.860 2.820 2.020 ;
        RECT  2.540 1.840 2.820 2.040 ;
        RECT  0.140 0.380 0.340 2.080 ;
        RECT  2.100 1.000 2.320 1.320 ;
        RECT  2.100 1.120 3.460 1.320 ;
        RECT  3.300 0.480 3.460 1.760 ;
        RECT  4.260 0.300 5.380 0.460 ;
        RECT  1.780 0.620 2.260 0.780 ;
        RECT  3.620 0.980 4.420 1.180 ;
        RECT  1.780 0.620 1.940 1.660 ;
        RECT  1.780 1.500 3.140 1.660 ;
        RECT  4.980 1.520 6.100 1.680 ;
        RECT  5.780 1.520 6.100 1.740 ;
        RECT  2.980 1.500 3.140 2.080 ;
        RECT  4.260 0.300 4.420 2.080 ;
        RECT  3.620 0.980 3.780 2.080 ;
        RECT  2.980 1.920 3.780 2.080 ;
        RECT  4.980 1.520 5.140 2.080 ;
        RECT  4.260 1.920 5.140 2.080 ;
        RECT  4.580 0.620 4.900 0.900 ;
        RECT  6.140 0.620 6.460 0.900 ;
        RECT  4.580 0.740 6.460 0.900 ;
        RECT  4.580 0.620 4.820 1.760 ;
        RECT  6.660 0.620 6.960 1.220 ;
        RECT  5.060 1.060 6.960 1.220 ;
        RECT  5.060 1.060 5.350 1.320 ;
        RECT  6.740 0.620 6.960 1.780 ;
        RECT  5.620 0.300 7.280 0.460 ;
        RECT  5.620 0.300 5.960 0.580 ;
        RECT  7.120 1.040 7.700 1.240 ;
        RECT  5.300 1.860 5.580 2.100 ;
        RECT  7.120 0.300 7.280 2.100 ;
        RECT  5.300 1.940 7.280 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END XNR3M4HM

MACRO XNR3M2HM
    CLASS CORE ;
    FOREIGN XNR3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        ANTENNAGATEAREA 0.136  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.684  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        ANTENNAGATEAREA 0.174  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.929  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 0.680 3.100 0.880 ;
        LAYER ME2 ;
        RECT  2.900 0.440 3.100 1.160 ;
        LAYER ME1 ;
        RECT  2.530 0.620 3.180 0.950 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.060 1.240 8.300 1.560 ;
        RECT  8.060 0.480 8.290 1.560 ;
        RECT  8.060 0.480 8.280 2.100 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        ANTENNAGATEAREA 0.156  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.367  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.430 1.440 6.630 1.640 ;
        LAYER ME2 ;
        RECT  6.360 1.240 6.700 1.960 ;
        LAYER ME1 ;
        RECT  6.380 1.380 6.690 1.780 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.560 1.430 7.720 2.540 ;
        RECT  3.980 1.440 4.140 2.540 ;
        RECT  0.660 1.800 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.560 -0.140 7.720 0.800 ;
        RECT  3.920 -0.140 4.120 0.820 ;
        RECT  0.620 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.380 0.620 1.660 1.700 ;
        RECT  1.060 0.300 2.940 0.460 ;
        RECT  0.140 1.480 1.220 1.640 ;
        RECT  1.060 0.300 1.220 2.020 ;
        RECT  1.060 1.860 2.860 2.020 ;
        RECT  2.580 1.840 2.860 2.040 ;
        RECT  0.140 0.380 0.340 2.080 ;
        RECT  2.140 1.000 2.360 1.320 ;
        RECT  2.140 1.120 3.500 1.320 ;
        RECT  3.340 0.480 3.500 1.760 ;
        RECT  4.300 0.300 5.420 0.460 ;
        RECT  1.820 0.620 2.300 0.780 ;
        RECT  3.660 0.980 4.460 1.180 ;
        RECT  1.820 0.620 1.980 1.660 ;
        RECT  1.820 1.500 3.180 1.660 ;
        RECT  5.020 1.520 6.220 1.680 ;
        RECT  5.900 1.520 6.220 1.740 ;
        RECT  3.020 1.500 3.180 2.080 ;
        RECT  4.300 0.300 4.460 2.080 ;
        RECT  3.660 0.980 3.820 2.080 ;
        RECT  3.020 1.920 3.820 2.080 ;
        RECT  5.020 1.520 5.180 2.080 ;
        RECT  4.300 1.920 5.180 2.080 ;
        RECT  4.620 0.620 4.940 0.900 ;
        RECT  6.260 0.620 6.580 0.900 ;
        RECT  4.620 0.740 6.580 0.900 ;
        RECT  4.620 0.620 4.860 1.760 ;
        RECT  6.780 0.620 7.080 1.220 ;
        RECT  5.100 1.060 7.080 1.220 ;
        RECT  5.100 1.060 5.390 1.320 ;
        RECT  6.860 0.620 7.080 1.780 ;
        RECT  5.660 0.300 7.400 0.460 ;
        RECT  5.660 0.300 6.000 0.580 ;
        RECT  7.240 1.040 7.820 1.240 ;
        RECT  5.340 1.860 5.620 2.100 ;
        RECT  7.240 0.300 7.400 2.100 ;
        RECT  5.340 1.940 7.400 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END XNR3M2HM

MACRO XNR3M1HM
    CLASS CORE ;
    FOREIGN XNR3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.655  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER ME1  ;
        ANTENNAGATEAREA 0.132  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.861  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 0.680 3.100 0.880 ;
        LAYER ME2 ;
        RECT  2.900 0.440 3.100 1.160 ;
        LAYER ME1 ;
        RECT  2.530 0.620 3.180 0.950 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.060 1.240 8.300 1.560 ;
        RECT  8.060 0.480 8.290 1.560 ;
        RECT  8.060 0.480 8.280 1.760 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.652  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.430 1.440 6.630 1.640 ;
        LAYER ME2 ;
        RECT  6.360 1.240 6.700 1.960 ;
        LAYER ME1 ;
        RECT  6.380 1.380 6.690 1.780 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.560 1.430 7.720 2.540 ;
        RECT  3.980 1.440 4.140 2.540 ;
        RECT  0.660 1.800 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.560 -0.140 7.720 0.800 ;
        RECT  3.920 -0.140 4.120 0.820 ;
        RECT  0.620 -0.140 0.860 0.760 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.380 0.620 1.660 1.700 ;
        RECT  1.060 0.300 2.940 0.460 ;
        RECT  0.140 1.480 1.220 1.640 ;
        RECT  1.060 0.300 1.220 2.020 ;
        RECT  1.060 1.860 2.860 2.020 ;
        RECT  2.580 1.840 2.860 2.040 ;
        RECT  0.140 0.470 0.340 2.080 ;
        RECT  2.140 1.000 2.360 1.320 ;
        RECT  2.140 1.120 3.500 1.320 ;
        RECT  3.340 0.470 3.500 1.760 ;
        RECT  4.300 0.300 5.420 0.460 ;
        RECT  1.820 0.620 2.300 0.780 ;
        RECT  3.660 0.980 4.460 1.180 ;
        RECT  1.820 0.620 1.980 1.660 ;
        RECT  1.820 1.500 3.180 1.660 ;
        RECT  5.020 1.520 6.220 1.680 ;
        RECT  5.900 1.520 6.220 1.740 ;
        RECT  3.020 1.500 3.180 2.080 ;
        RECT  4.300 0.300 4.460 2.080 ;
        RECT  3.660 0.980 3.820 2.080 ;
        RECT  3.020 1.920 3.820 2.080 ;
        RECT  5.020 1.520 5.180 2.080 ;
        RECT  4.300 1.920 5.180 2.080 ;
        RECT  4.620 0.620 4.940 0.900 ;
        RECT  6.260 0.620 6.580 0.900 ;
        RECT  4.620 0.740 6.580 0.900 ;
        RECT  4.620 0.620 4.860 1.760 ;
        RECT  6.780 0.620 7.080 1.220 ;
        RECT  5.100 1.060 7.080 1.220 ;
        RECT  5.100 1.060 5.390 1.320 ;
        RECT  6.860 0.620 7.080 1.780 ;
        RECT  5.660 0.300 7.400 0.460 ;
        RECT  5.660 0.300 6.000 0.550 ;
        RECT  7.240 1.040 7.820 1.240 ;
        RECT  5.340 1.860 5.620 2.100 ;
        RECT  7.240 0.300 7.400 2.100 ;
        RECT  5.340 1.940 7.400 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END XNR3M1HM

MACRO XNR3M0HM
    CLASS CORE ;
    FOREIGN XNR3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.740  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER ME1  ;
        ANTENNAGATEAREA 0.132  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.861  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 0.680 3.100 0.880 ;
        LAYER ME2 ;
        RECT  2.900 0.440 3.100 1.160 ;
        LAYER ME1 ;
        RECT  2.530 0.620 3.180 0.950 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.060 1.240 8.300 1.560 ;
        RECT  8.060 0.530 8.290 1.560 ;
        RECT  8.060 0.530 8.280 1.760 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER ME1  ;
        ANTENNAGATEAREA 0.132  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.797  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.430 1.440 6.630 1.640 ;
        LAYER ME2 ;
        RECT  6.360 1.240 6.700 1.960 ;
        LAYER ME1 ;
        RECT  6.380 1.380 6.690 1.780 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.560 1.430 7.720 2.540 ;
        RECT  3.980 1.440 4.140 2.540 ;
        RECT  0.660 1.800 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.560 -0.140 7.720 0.850 ;
        RECT  3.920 -0.140 4.120 0.820 ;
        RECT  0.620 -0.140 0.860 0.750 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.380 0.620 1.660 1.700 ;
        RECT  1.060 0.300 2.940 0.460 ;
        RECT  0.140 1.480 1.220 1.640 ;
        RECT  1.060 0.300 1.220 2.020 ;
        RECT  1.060 1.860 2.860 2.020 ;
        RECT  2.580 1.840 2.860 2.040 ;
        RECT  0.140 0.470 0.340 2.080 ;
        RECT  2.140 1.000 2.360 1.320 ;
        RECT  2.140 1.120 3.500 1.320 ;
        RECT  3.340 0.470 3.500 1.760 ;
        RECT  4.300 0.300 5.420 0.460 ;
        RECT  1.820 0.620 2.300 0.780 ;
        RECT  3.660 0.980 4.460 1.180 ;
        RECT  1.820 0.620 1.980 1.660 ;
        RECT  1.820 1.500 3.180 1.660 ;
        RECT  5.020 1.520 6.220 1.680 ;
        RECT  5.900 1.520 6.220 1.740 ;
        RECT  3.020 1.500 3.180 2.080 ;
        RECT  4.300 0.300 4.460 2.080 ;
        RECT  3.660 0.980 3.820 2.080 ;
        RECT  3.020 1.920 3.820 2.080 ;
        RECT  5.020 1.520 5.180 2.080 ;
        RECT  4.300 1.920 5.180 2.080 ;
        RECT  4.620 0.620 4.940 0.900 ;
        RECT  6.260 0.620 6.580 0.900 ;
        RECT  4.620 0.740 6.580 0.900 ;
        RECT  4.620 0.620 4.860 1.760 ;
        RECT  6.780 0.620 7.080 1.220 ;
        RECT  5.100 1.060 7.080 1.220 ;
        RECT  5.100 1.060 5.390 1.320 ;
        RECT  6.860 0.620 7.080 1.780 ;
        RECT  5.660 0.300 7.400 0.460 ;
        RECT  5.660 0.300 6.000 0.550 ;
        RECT  7.240 1.040 7.820 1.240 ;
        RECT  5.340 1.860 5.620 2.100 ;
        RECT  7.240 0.300 7.400 2.100 ;
        RECT  5.340 1.940 7.400 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END XNR3M0HM

MACRO XNR2M4HM
    CLASS CORE ;
    FOREIGN XNR2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.446  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.176  LAYER ME1  ;
        ANTENNAGATEAREA 0.176  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.095  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 0.680 3.100 0.880 ;
        LAYER ME2 ;
        RECT  2.900 0.440 3.100 1.160 ;
        LAYER ME1 ;
        RECT  2.490 0.620 3.140 1.020 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.740 1.240 5.100 1.560 ;
        RECT  4.740 0.430 4.970 1.560 ;
        RECT  4.740 0.430 4.960 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.260 1.470 5.460 2.540 ;
        RECT  4.240 1.430 4.400 2.540 ;
        RECT  0.660 1.800 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.260 -0.140 5.460 0.710 ;
        RECT  4.240 -0.140 4.400 0.750 ;
        RECT  0.660 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.620 1.620 1.700 ;
        RECT  1.020 0.300 3.220 0.460 ;
        RECT  0.140 1.480 1.180 1.640 ;
        RECT  1.020 0.300 1.180 2.020 ;
        RECT  1.020 1.860 3.110 2.020 ;
        RECT  2.830 1.840 3.110 2.040 ;
        RECT  0.140 0.380 0.340 2.080 ;
        RECT  2.100 1.000 2.320 1.340 ;
        RECT  2.100 1.180 3.760 1.340 ;
        RECT  3.600 0.480 3.760 1.760 ;
        RECT  1.780 0.620 2.260 0.780 ;
        RECT  3.920 1.040 4.520 1.240 ;
        RECT  1.780 0.620 1.940 1.660 ;
        RECT  1.780 1.500 3.430 1.660 ;
        RECT  3.270 1.500 3.430 2.080 ;
        RECT  3.920 1.040 4.080 2.080 ;
        RECT  3.270 1.920 4.080 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END XNR2M4HM

MACRO XNR2M2HM
    CLASS CORE ;
    FOREIGN XNR2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.571  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.216  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 1.240 4.300 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.681  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.340 3.280 0.540 ;
        RECT  2.980 1.170 3.260 1.660 ;
        RECT  2.860 0.340 3.020 1.330 ;
        RECT  1.900 1.170 3.260 1.330 ;
        RECT  1.900 1.170 2.300 1.760 ;
        RECT  1.900 0.620 2.220 1.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.790 4.300 2.540 ;
        RECT  0.680 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.020 -0.140 4.300 0.770 ;
        RECT  0.660 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.620 1.620 1.760 ;
        RECT  1.020 0.300 2.700 0.460 ;
        RECT  2.470 0.300 2.700 0.630 ;
        RECT  0.140 1.480 1.180 1.640 ;
        RECT  1.020 0.300 1.180 2.100 ;
        RECT  0.140 0.400 0.340 2.080 ;
        RECT  2.460 1.520 2.740 2.100 ;
        RECT  1.020 1.940 2.740 2.100 ;
        RECT  3.180 0.700 3.740 0.980 ;
        RECT  3.540 0.490 3.740 2.100 ;
        RECT  3.120 1.880 3.740 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END XNR2M2HM

MACRO XNR2M1HM
    CLASS CORE ;
    FOREIGN XNR2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        ANTENNAGATEAREA 0.104  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.487  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.010 0.700 1.210 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.950 0.860 1.290 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.188  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 1.220 4.300 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.597  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.340 3.280 0.540 ;
        RECT  2.980 1.170 3.260 1.680 ;
        RECT  2.860 0.340 3.020 1.330 ;
        RECT  1.900 1.170 3.260 1.330 ;
        RECT  1.900 1.170 2.300 1.680 ;
        RECT  1.900 0.620 2.180 1.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.060 1.790 4.260 2.540 ;
        RECT  0.680 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.770 ;
        RECT  0.660 -0.140 0.860 0.770 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.620 1.620 1.680 ;
        RECT  1.020 0.300 2.700 0.460 ;
        RECT  2.470 0.300 2.700 0.630 ;
        RECT  0.140 1.480 1.180 1.640 ;
        RECT  1.020 0.300 1.180 2.100 ;
        RECT  0.140 0.490 0.340 2.080 ;
        RECT  2.460 1.520 2.740 2.100 ;
        RECT  1.020 1.940 2.740 2.100 ;
        RECT  3.180 0.700 3.740 0.980 ;
        RECT  3.540 0.490 3.740 2.100 ;
        RECT  3.120 1.900 3.740 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END XNR2M1HM

MACRO XNR2M0HM
    CLASS CORE ;
    FOREIGN XNR2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.387  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.840 2.300 1.160 ;
        RECT  1.900 0.620 2.180 1.680 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.395  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.570 1.050 0.770 1.250 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.770 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.970 0.860 1.320 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.500 1.220 3.900 1.560 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.660 1.790 3.860 2.540 ;
        RECT  0.680 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.660 -0.140 3.860 0.560 ;
        RECT  0.660 -0.140 0.860 0.810 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.620 1.620 1.680 ;
        RECT  1.020 0.300 2.760 0.460 ;
        RECT  2.470 0.300 2.760 0.520 ;
        RECT  0.140 1.480 1.180 1.640 ;
        RECT  2.340 1.520 2.740 1.740 ;
        RECT  1.020 0.300 1.180 2.100 ;
        RECT  0.140 0.520 0.340 2.080 ;
        RECT  2.340 1.520 2.500 2.100 ;
        RECT  1.020 1.940 2.500 2.100 ;
        RECT  3.100 0.340 3.380 0.590 ;
        RECT  3.100 0.340 3.340 0.980 ;
        RECT  2.720 0.760 3.340 0.980 ;
        RECT  3.140 0.340 3.340 2.100 ;
        RECT  2.720 1.900 3.340 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END XNR2M0HM

MACRO WTBP2HM
    CLASS CORE ;
    FOREIGN WTBP2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VBP
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.470 0.540 2.100 ;
        END
    END VBP
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.800 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.800 0.140 ;
        RECT  0.300 -0.140 0.500 0.830 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.800 1.140 ;
    END
END WTBP2HM

MACRO WTBN2HM
    CLASS CORE ;
    FOREIGN WTBN2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VBN
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.440 0.500 0.830 ;
        END
    END VBN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.800 2.540 ;
        RECT  0.300 1.470 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.800 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.800 1.140 ;
    END
END WTBN2HM

MACRO WTBB2HM
    CLASS CORE ;
    FOREIGN WTBB2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VBN
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.440 0.500 0.830 ;
        END
    END VBN
    PIN VBP
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.470 0.540 2.100 ;
        END
    END VBP
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.800 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.800 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.800 1.140 ;
    END
END WTBB2HM

MACRO WT2HM
    CLASS CORE ;
    FOREIGN WT2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.800 2.540 ;
        RECT  0.300 1.510 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.800 0.140 ;
        RECT  0.300 -0.140 0.500 0.830 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.800 1.140 ;
    END
END WT2HM

MACRO TIE1HM
    CLASS CORE ;
    FOREIGN TIE1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.231  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.520 1.100 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.240 1.480 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.760 -0.140 0.960 0.760 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 0.480 0.440 1.210 ;
        RECT  0.240 1.010 0.660 1.210 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END TIE1HM

MACRO TIE0HM
    CLASS CORE ;
    FOREIGN TIE0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.190  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.430 1.100 1.160 ;
        RECT  0.720 0.430 1.100 0.630 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.760 1.640 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.240 -0.140 0.440 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 1.220 0.660 1.420 ;
        RECT  0.240 1.220 0.440 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END TIE0HM

MACRO SDFZRM8HM
    CLASS CORE ;
    FOREIGN SDFZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        ANTENNAGATEAREA 0.146  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.628  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.312  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.320 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.190  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.300 0.430 16.500 1.720 ;
        RECT  14.940 0.900 16.500 1.100 ;
        RECT  15.100 0.430 15.300 1.100 ;
        RECT  14.940 0.900 15.140 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  18.540 0.430 18.740 2.100 ;
        RECT  17.500 1.420 18.740 1.630 ;
        RECT  18.500 0.660 18.740 1.630 ;
        RECT  17.500 0.660 18.740 0.860 ;
        RECT  17.500 1.420 17.700 2.100 ;
        RECT  17.500 0.430 17.700 0.860 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.570 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 19.600 2.540 ;
        RECT  19.060 1.460 19.260 2.540 ;
        RECT  18.020 1.840 18.220 2.540 ;
        RECT  16.980 1.480 17.180 2.540 ;
        RECT  15.620 1.840 15.820 2.540 ;
        RECT  14.260 1.840 14.460 2.540 ;
        RECT  12.980 1.840 13.260 2.540 ;
        RECT  10.600 1.800 10.760 2.540 ;
        RECT  9.160 2.080 9.440 2.540 ;
        RECT  5.820 1.840 6.020 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 19.600 0.140 ;
        RECT  19.060 -0.140 19.260 0.710 ;
        RECT  17.980 -0.140 18.260 0.500 ;
        RECT  16.950 -0.140 17.150 0.710 ;
        RECT  15.620 -0.140 15.820 0.710 ;
        RECT  14.580 -0.140 14.780 0.710 ;
        RECT  13.600 -0.140 13.760 0.700 ;
        RECT  10.600 -0.140 10.880 0.500 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.380 1.420 0.580 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.380 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.340 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  6.780 0.620 7.060 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.500 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.300 0.300 7.500 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  8.040 0.620 8.240 1.080 ;
        RECT  8.040 0.880 9.620 1.080 ;
        RECT  8.040 0.620 8.220 1.740 ;
        RECT  8.040 1.540 8.420 1.740 ;
        RECT  8.880 1.240 9.080 1.600 ;
        RECT  9.840 0.620 10.120 1.600 ;
        RECT  8.880 1.440 10.120 1.600 ;
        RECT  9.920 0.620 10.120 1.780 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.340 0.960 ;
        RECT  10.280 1.360 10.920 1.560 ;
        RECT  5.300 1.480 6.340 1.680 ;
        RECT  5.300 1.480 5.500 1.920 ;
        RECT  8.840 1.760 9.760 1.920 ;
        RECT  6.180 0.800 6.340 2.100 ;
        RECT  9.600 1.760 9.760 2.100 ;
        RECT  8.840 1.760 9.000 2.100 ;
        RECT  6.180 1.940 9.000 2.100 ;
        RECT  10.280 1.360 10.440 2.100 ;
        RECT  9.600 1.940 10.440 2.100 ;
        RECT  11.040 0.300 11.540 0.600 ;
        RECT  7.680 0.300 8.560 0.460 ;
        RECT  9.360 0.300 10.440 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  9.360 0.300 9.520 0.720 ;
        RECT  8.400 0.560 9.520 0.720 ;
        RECT  10.280 0.300 10.440 0.940 ;
        RECT  10.280 0.780 11.600 0.940 ;
        RECT  11.380 0.780 11.600 1.100 ;
        RECT  7.680 0.300 7.880 1.540 ;
        RECT  11.760 0.300 11.960 1.700 ;
        RECT  11.480 1.540 11.960 1.700 ;
        RECT  12.660 0.620 13.120 0.900 ;
        RECT  12.300 0.300 13.440 0.460 ;
        RECT  12.300 0.300 12.500 0.700 ;
        RECT  13.280 0.300 13.440 1.280 ;
        RECT  12.120 1.080 13.840 1.280 ;
        RECT  12.120 1.080 12.280 2.020 ;
        RECT  10.980 1.860 12.280 2.020 ;
        RECT  16.660 1.020 17.920 1.220 ;
        RECT  14.100 0.430 14.300 1.680 ;
        RECT  12.760 1.480 14.780 1.680 ;
        RECT  15.300 1.520 16.140 1.680 ;
        RECT  14.620 1.480 14.780 2.100 ;
        RECT  15.980 1.520 16.140 2.100 ;
        RECT  15.300 1.520 15.460 2.100 ;
        RECT  14.620 1.940 15.460 2.100 ;
        RECT  16.660 1.020 16.820 2.100 ;
        RECT  15.980 1.940 16.820 2.100 ;
        LAYER VI1 ;
        RECT  6.780 1.200 6.980 1.400 ;
        RECT  7.680 1.200 7.880 1.400 ;
        RECT  9.920 0.960 10.120 1.160 ;
        RECT  10.620 1.360 10.820 1.560 ;
        RECT  11.140 0.400 11.340 0.600 ;
        RECT  11.760 0.960 11.960 1.160 ;
        RECT  12.300 0.400 12.500 0.600 ;
        RECT  12.820 0.620 13.020 0.820 ;
        LAYER ME2 ;
        RECT  6.680 1.200 7.980 1.400 ;
        RECT  9.840 0.960 12.020 1.160 ;
        RECT  11.040 0.400 12.600 0.600 ;
        RECT  12.820 0.520 13.020 1.560 ;
        RECT  10.520 1.360 13.020 1.560 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  10.810 1.090 12.520 2.400 ;
        RECT  0.000 1.140 7.770 2.400 ;
        RECT  8.800 1.140 19.600 2.400 ;
        RECT  0.000 1.200 19.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 19.600 1.080 ;
        RECT  4.080 0.000 19.600 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 10.810 1.140 ;
        RECT  12.520 0.000 19.600 1.140 ;
        RECT  7.770 0.000 8.800 1.200 ;
    END
END SDFZRM8HM

MACRO SDFZRM4HM
    CLASS CORE ;
    FOREIGN SDFZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        ANTENNAGATEAREA 0.078  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.933  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.312  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.380 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.200 0.900 13.760 1.100 ;
        RECT  13.560 0.390 13.760 1.100 ;
        RECT  13.400 0.900 13.600 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.600 1.420 15.500 1.630 ;
        RECT  15.300 0.660 15.500 1.630 ;
        RECT  14.600 0.660 15.500 0.860 ;
        RECT  14.600 1.420 14.800 2.100 ;
        RECT  14.600 0.430 14.800 0.860 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.570 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  15.120 1.840 15.320 2.540 ;
        RECT  14.080 1.840 14.280 2.540 ;
        RECT  12.720 1.840 12.920 2.540 ;
        RECT  11.630 1.840 11.910 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.820 1.840 6.020 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  15.080 -0.140 15.360 0.500 ;
        RECT  14.080 -0.140 14.280 0.670 ;
        RECT  13.040 -0.140 13.240 0.670 ;
        RECT  12.060 -0.140 12.220 0.700 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.380 1.420 0.580 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.380 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.340 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  6.780 0.620 7.060 1.400 ;
        RECT  6.540 1.220 7.060 1.400 ;
        RECT  6.540 1.220 6.740 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.480 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.220 0.300 7.480 0.660 ;
        RECT  7.220 0.300 7.380 1.780 ;
        RECT  6.980 1.580 7.380 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  7.960 0.880 9.460 1.080 ;
        RECT  7.960 0.620 8.160 1.780 ;
        RECT  7.880 1.580 8.160 1.780 ;
        RECT  7.640 0.300 8.560 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  8.400 0.560 9.880 0.720 ;
        RECT  7.640 0.300 7.800 1.000 ;
        RECT  9.720 0.560 9.880 1.090 ;
        RECT  7.540 0.850 7.700 1.490 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.340 0.960 ;
        RECT  5.300 1.500 6.340 1.680 ;
        RECT  8.420 1.720 9.560 1.920 ;
        RECT  6.180 0.800 6.340 2.100 ;
        RECT  5.300 1.500 5.500 2.050 ;
        RECT  8.420 1.720 8.580 2.100 ;
        RECT  6.180 1.940 8.580 2.100 ;
        RECT  9.400 1.900 10.080 2.100 ;
        RECT  10.040 0.300 10.200 1.460 ;
        RECT  8.700 1.300 10.200 1.460 ;
        RECT  9.720 1.300 9.920 1.720 ;
        RECT  11.120 0.620 11.580 0.900 ;
        RECT  10.560 0.300 11.900 0.460 ;
        RECT  10.560 0.300 10.760 0.660 ;
        RECT  11.740 0.300 11.900 1.280 ;
        RECT  10.580 1.080 12.300 1.280 ;
        RECT  10.580 1.080 10.740 1.950 ;
        RECT  13.920 1.020 15.020 1.220 ;
        RECT  12.560 0.390 12.760 1.680 ;
        RECT  11.220 1.480 13.240 1.680 ;
        RECT  13.920 1.020 14.080 1.680 ;
        RECT  13.080 1.480 13.240 2.100 ;
        RECT  13.760 1.520 13.920 2.100 ;
        RECT  13.080 1.940 13.920 2.100 ;
        LAYER VI1 ;
        RECT  9.200 1.720 9.400 1.920 ;
        RECT  11.280 0.620 11.480 0.820 ;
        LAYER ME2 ;
        RECT  11.280 0.520 11.480 1.920 ;
        RECT  9.100 1.720 11.480 1.920 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  8.800 1.090 10.980 2.400 ;
        RECT  0.000 1.140 5.840 2.400 ;
        RECT  8.800 1.140 15.600 2.400 ;
        RECT  0.000 1.200 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.080 ;
        RECT  4.080 0.000 15.600 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 8.800 1.140 ;
        RECT  10.980 0.000 15.600 1.140 ;
        RECT  5.840 0.000 8.800 1.200 ;
    END
END SDFZRM4HM

MACRO SDFZRM2HM
    CLASS CORE ;
    FOREIGN SDFZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        ANTENNAGATEAREA 0.078  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.933  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.312  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.320 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.900 0.390 13.100 1.160 ;
        RECT  12.740 0.950 12.940 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.900 1.440 14.300 2.100 ;
        RECT  14.100 0.470 14.300 2.100 ;
        RECT  13.900 0.470 14.300 0.670 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.570 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.400 2.540 ;
        RECT  13.420 1.840 13.620 2.540 ;
        RECT  11.640 1.840 11.840 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.820 1.840 6.020 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.400 0.140 ;
        RECT  13.420 -0.140 13.620 0.670 ;
        RECT  11.780 -0.140 11.940 0.610 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.380 1.420 0.580 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.380 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.340 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  6.780 0.620 7.060 1.400 ;
        RECT  6.540 1.220 7.060 1.400 ;
        RECT  6.540 1.220 6.740 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.480 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.220 0.300 7.480 0.660 ;
        RECT  7.220 0.300 7.380 1.780 ;
        RECT  6.980 1.580 7.380 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  7.960 0.880 9.460 1.080 ;
        RECT  7.960 0.620 8.160 1.780 ;
        RECT  7.880 1.580 8.160 1.780 ;
        RECT  7.640 0.300 8.560 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  8.400 0.560 9.880 0.720 ;
        RECT  7.640 0.300 7.800 1.000 ;
        RECT  9.720 0.560 9.880 1.090 ;
        RECT  7.540 0.850 7.700 1.490 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.340 0.960 ;
        RECT  5.300 1.500 6.340 1.680 ;
        RECT  8.420 1.720 9.560 1.920 ;
        RECT  6.180 0.800 6.340 2.100 ;
        RECT  5.300 1.500 5.500 2.050 ;
        RECT  8.420 1.720 8.580 2.100 ;
        RECT  6.180 1.940 8.580 2.100 ;
        RECT  9.400 1.900 10.080 2.100 ;
        RECT  10.040 0.300 10.200 1.460 ;
        RECT  8.700 1.300 10.200 1.460 ;
        RECT  9.720 1.300 9.920 1.720 ;
        RECT  10.920 0.620 11.380 0.900 ;
        RECT  12.060 1.000 12.260 1.280 ;
        RECT  10.560 1.080 12.260 1.280 ;
        RECT  10.560 0.380 10.760 2.070 ;
        RECT  12.320 0.300 12.580 0.580 ;
        RECT  11.220 1.480 12.580 1.680 ;
        RECT  13.580 0.940 13.740 1.680 ;
        RECT  13.100 1.520 13.740 1.680 ;
        RECT  12.420 0.300 12.580 2.100 ;
        RECT  13.100 1.520 13.260 2.100 ;
        RECT  12.420 1.940 13.260 2.100 ;
        LAYER VI1 ;
        RECT  9.200 1.720 9.400 1.920 ;
        RECT  11.080 0.620 11.280 0.820 ;
        LAYER ME2 ;
        RECT  11.080 0.520 11.280 1.920 ;
        RECT  9.100 1.720 11.280 1.920 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  8.800 1.090 10.980 2.400 ;
        RECT  0.000 1.140 5.840 2.400 ;
        RECT  8.800 1.140 14.400 2.400 ;
        RECT  0.000 1.200 14.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.400 1.080 ;
        RECT  4.080 0.000 14.400 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 8.800 1.140 ;
        RECT  10.980 0.000 14.400 1.140 ;
        RECT  5.840 0.000 8.800 1.200 ;
    END
END SDFZRM2HM

MACRO SDFZRM1HM
    CLASS CORE ;
    FOREIGN SDFZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        ANTENNAGATEAREA 0.053  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.288  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        ANTENNAGATEAREA 0.065  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.099  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.320 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.354  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.900 0.390 13.100 1.160 ;
        RECT  12.740 0.950 12.940 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.900 1.800 14.300 2.000 ;
        RECT  14.100 0.390 14.300 2.000 ;
        RECT  13.900 0.390 14.300 0.590 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.600 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.400 2.540 ;
        RECT  13.420 1.840 13.620 2.540 ;
        RECT  11.640 1.840 11.840 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.900 1.840 6.100 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.400 0.140 ;
        RECT  13.420 -0.140 13.620 0.670 ;
        RECT  11.780 -0.140 11.940 0.610 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.400 1.420 0.600 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.400 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.320 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  1.880 1.760 2.080 2.100 ;
        RECT  6.780 0.620 7.060 1.400 ;
        RECT  6.580 1.220 6.780 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.480 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.220 0.300 7.480 0.660 ;
        RECT  7.220 0.300 7.380 1.780 ;
        RECT  7.020 1.580 7.380 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  7.960 0.880 9.460 1.080 ;
        RECT  7.960 0.620 8.160 1.780 ;
        RECT  7.880 1.580 8.160 1.780 ;
        RECT  7.640 0.300 8.560 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  8.400 0.560 9.880 0.720 ;
        RECT  7.640 0.300 7.800 1.000 ;
        RECT  9.720 0.560 9.880 1.090 ;
        RECT  7.540 0.850 7.700 1.490 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.420 0.960 ;
        RECT  5.300 1.500 6.420 1.680 ;
        RECT  8.420 1.720 9.560 1.920 ;
        RECT  6.260 0.800 6.420 2.100 ;
        RECT  5.300 1.500 5.500 2.100 ;
        RECT  8.420 1.720 8.580 2.100 ;
        RECT  6.260 1.940 8.580 2.100 ;
        RECT  9.400 1.900 10.080 2.100 ;
        RECT  10.040 0.300 10.200 1.460 ;
        RECT  8.700 1.300 10.200 1.460 ;
        RECT  9.720 1.300 9.920 1.720 ;
        RECT  10.920 0.620 11.380 0.900 ;
        RECT  12.060 1.000 12.260 1.280 ;
        RECT  10.560 1.080 12.260 1.280 ;
        RECT  10.560 0.380 10.760 2.070 ;
        RECT  12.320 0.300 12.580 0.580 ;
        RECT  11.220 1.480 12.580 1.680 ;
        RECT  13.580 0.940 13.740 1.680 ;
        RECT  13.100 1.520 13.740 1.680 ;
        RECT  12.420 0.300 12.580 2.100 ;
        RECT  13.100 1.520 13.260 2.100 ;
        RECT  12.420 1.940 13.260 2.100 ;
        LAYER VI1 ;
        RECT  9.200 1.720 9.400 1.920 ;
        RECT  11.080 0.620 11.280 0.820 ;
        LAYER ME2 ;
        RECT  11.080 0.520 11.280 1.920 ;
        RECT  9.100 1.720 11.280 1.920 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  8.800 1.090 10.980 2.400 ;
        RECT  0.000 1.140 5.840 2.400 ;
        RECT  8.800 1.140 14.400 2.400 ;
        RECT  0.000 1.200 14.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.400 1.080 ;
        RECT  4.080 0.000 14.400 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 8.800 1.140 ;
        RECT  10.980 0.000 14.400 1.140 ;
        RECT  5.840 0.000 8.800 1.200 ;
    END
END SDFZRM1HM

MACRO SDFSM8HM
    CLASS CORE ;
    FOREIGN SDFSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.180 0.840 7.500 1.160 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.620 3.240 3.100 3.720 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.960  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.440 1.900 2.080 ;
        RECT  0.900 0.660 1.900 0.860 ;
        RECT  1.700 0.440 1.900 0.860 ;
        RECT  0.660 1.440 1.900 1.640 ;
        RECT  0.900 0.660 1.100 1.640 ;
        RECT  0.660 0.660 1.900 0.830 ;
        RECT  0.660 1.440 0.860 2.080 ;
        RECT  0.660 0.440 0.860 0.830 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.116  LAYER ME1  ;
        ANTENNADIFFAREA 1.027  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.900 1.860 8.300 2.060 ;
        RECT  8.100 0.420 8.300 2.060 ;
        RECT  7.900 0.420 8.300 0.620 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.242  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.960 1.120 4.360 1.500 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.061  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 3.550 1.160 4.000 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.550 0.700 4.100 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.460 1.500 8.660 3.300 ;
        RECT  7.380 2.260 7.580 3.300 ;
        RECT  3.260 1.860 3.460 2.540 ;
        RECT  2.860 2.260 3.140 2.640 ;
        RECT  2.220 1.860 2.420 2.540 ;
        RECT  1.180 1.860 1.380 2.540 ;
        RECT  0.660 2.260 0.940 2.960 ;
        RECT  0.140 1.500 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.460 -0.140 8.660 0.660 ;
        RECT  7.380 -0.140 7.580 0.660 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.710 ;
        RECT  0.000 4.660 8.800 4.940 ;
        RECT  8.460 4.180 8.660 4.940 ;
        RECT  7.380 4.180 7.580 4.940 ;
        RECT  4.740 4.480 5.020 4.940 ;
        RECT  2.940 4.240 3.140 4.940 ;
        RECT  0.660 4.260 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.120 1.520 3.280 ;
        RECT  1.360 3.120 1.520 3.870 ;
        RECT  1.360 3.670 2.000 3.870 ;
        RECT  0.140 3.030 0.340 4.290 ;
        RECT  2.180 3.120 2.460 4.160 ;
        RECT  2.740 0.440 2.940 0.860 ;
        RECT  2.220 0.660 2.940 0.860 ;
        RECT  1.480 1.040 2.420 1.240 ;
        RECT  2.220 0.660 2.420 1.570 ;
        RECT  3.480 1.060 3.680 1.570 ;
        RECT  2.220 1.380 3.680 1.570 ;
        RECT  2.740 1.380 2.940 2.080 ;
        RECT  3.980 3.780 4.640 4.000 ;
        RECT  3.980 3.780 4.260 4.160 ;
        RECT  3.280 3.440 5.140 3.600 ;
        RECT  3.280 3.440 3.480 3.760 ;
        RECT  4.860 3.360 5.140 4.000 ;
        RECT  4.860 3.840 6.020 4.000 ;
        RECT  5.740 3.840 6.020 4.160 ;
        RECT  1.660 2.720 2.660 2.880 ;
        RECT  3.280 2.720 6.060 2.880 ;
        RECT  2.500 2.800 3.420 2.960 ;
        RECT  1.660 2.720 1.860 3.020 ;
        RECT  3.660 0.320 6.260 0.480 ;
        RECT  3.660 0.320 3.820 0.860 ;
        RECT  3.100 0.660 3.820 0.860 ;
        RECT  6.060 0.320 6.260 0.880 ;
        RECT  3.100 0.660 3.260 1.220 ;
        RECT  2.700 1.060 3.260 1.220 ;
        RECT  4.880 0.320 5.040 1.620 ;
        RECT  4.880 1.460 5.860 1.620 ;
        RECT  5.580 1.460 5.860 1.760 ;
        RECT  5.380 0.660 5.740 0.820 ;
        RECT  5.580 0.660 5.740 1.200 ;
        RECT  5.580 1.040 6.180 1.200 ;
        RECT  6.020 1.040 6.180 1.760 ;
        RECT  6.020 1.600 6.490 1.760 ;
        RECT  2.620 3.920 3.460 4.080 ;
        RECT  1.660 4.140 1.860 4.480 ;
        RECT  3.300 3.920 3.460 4.480 ;
        RECT  4.420 4.160 5.340 4.320 ;
        RECT  2.620 3.920 2.780 4.480 ;
        RECT  1.660 4.320 2.780 4.480 ;
        RECT  3.300 4.320 4.580 4.480 ;
        RECT  6.340 4.050 6.540 4.480 ;
        RECT  5.180 4.320 6.540 4.480 ;
        RECT  6.220 2.700 6.660 2.860 ;
        RECT  4.360 3.040 6.380 3.200 ;
        RECT  6.220 2.700 6.380 3.200 ;
        RECT  3.380 3.120 4.640 3.280 ;
        RECT  5.320 3.480 7.020 3.640 ;
        RECT  6.820 3.080 7.020 4.330 ;
        RECT  6.400 1.030 7.020 1.230 ;
        RECT  6.820 0.380 7.020 1.760 ;
        RECT  4.130 0.640 4.680 0.800 ;
        RECT  7.780 0.980 7.940 1.700 ;
        RECT  7.350 1.540 7.940 1.700 ;
        RECT  4.520 0.640 4.680 2.080 ;
        RECT  3.820 1.690 4.020 2.080 ;
        RECT  4.520 1.780 5.100 2.080 ;
        RECT  7.350 1.540 7.510 2.080 ;
        RECT  3.820 1.920 7.510 2.080 ;
        RECT  7.940 2.720 8.140 4.350 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.550 3.640 ;
        RECT  0.000 1.180 8.800 3.640 ;
        RECT  0.000 1.140 1.970 3.660 ;
        RECT  6.450 1.140 8.800 3.660 ;
        RECT  6.320 1.180 8.800 3.660 ;
        RECT  4.560 1.180 5.440 3.880 ;
        LAYER VTNH ;
        RECT  5.440 3.640 6.320 4.800 ;
        RECT  1.970 3.640 4.560 4.800 ;
        RECT  0.000 3.660 4.560 4.800 ;
        RECT  5.440 3.660 8.800 4.800 ;
        RECT  0.000 3.880 8.800 4.800 ;
        RECT  0.000 0.000 8.800 1.140 ;
        RECT  3.550 0.000 6.450 1.180 ;
    END
END SDFSM8HM

MACRO SDFSM4HM
    CLASS CORE ;
    FOREIGN SDFSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.190 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.400 0.440 14.700 0.800 ;
        RECT  14.400 0.440 14.560 1.760 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.540 1.440 16.300 1.640 ;
        RECT  16.100 0.740 16.300 1.640 ;
        RECT  15.540 0.740 16.300 0.900 ;
        RECT  15.540 1.440 15.740 2.080 ;
        RECT  15.540 0.450 15.740 0.900 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.250  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.740 1.430 12.620 1.590 ;
        RECT  12.100 1.120 12.620 1.590 ;
        RECT  10.120 1.940 10.900 2.100 ;
        RECT  10.740 1.430 10.900 2.100 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.400 2.540 ;
        RECT  16.060 1.840 16.260 2.540 ;
        RECT  15.040 1.440 15.200 2.540 ;
        RECT  13.760 1.800 13.920 2.540 ;
        RECT  12.100 2.080 12.380 2.540 ;
        RECT  11.060 1.840 11.260 2.540 ;
        RECT  8.020 2.080 8.300 2.540 ;
        RECT  4.360 2.020 4.560 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.400 0.140 ;
        RECT  16.060 -0.140 16.260 0.560 ;
        RECT  15.020 -0.140 15.220 0.650 ;
        RECT  13.700 -0.140 13.980 0.500 ;
        RECT  12.380 -0.140 12.660 0.320 ;
        RECT  10.980 -0.140 11.140 0.650 ;
        RECT  7.400 -0.140 7.600 0.560 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.300 ;
        RECT  3.700 1.100 4.820 1.300 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.700 4.880 1.860 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.720 1.700 4.880 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.700 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.520 1.740 5.720 2.100 ;
        RECT  4.720 1.940 5.720 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.640 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.640 5.460 1.510 ;
        RECT  5.040 1.350 5.460 1.510 ;
        RECT  5.040 1.350 5.240 1.780 ;
        RECT  6.460 0.900 7.880 1.060 ;
        RECT  7.680 0.900 7.880 1.220 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  6.040 1.240 6.660 1.400 ;
        RECT  6.040 1.240 6.240 2.020 ;
        RECT  8.040 0.350 8.580 0.550 ;
        RECT  6.920 1.240 7.120 1.600 ;
        RECT  8.040 0.350 8.200 1.600 ;
        RECT  6.920 1.440 8.980 1.600 ;
        RECT  8.780 1.440 8.980 1.780 ;
        RECT  9.140 0.980 9.480 1.180 ;
        RECT  6.400 1.760 8.620 1.920 ;
        RECT  8.460 1.760 8.620 2.100 ;
        RECT  6.400 1.760 6.680 2.100 ;
        RECT  9.140 0.980 9.300 2.100 ;
        RECT  8.460 1.940 9.300 2.100 ;
        RECT  8.760 0.660 9.900 0.820 ;
        RECT  8.760 0.660 8.960 1.200 ;
        RECT  9.740 0.660 9.900 1.270 ;
        RECT  8.860 0.300 10.220 0.500 ;
        RECT  10.060 0.300 10.220 1.760 ;
        RECT  9.460 1.480 10.220 1.760 ;
        RECT  11.620 0.620 11.900 0.960 ;
        RECT  11.620 0.800 12.940 0.960 ;
        RECT  12.780 1.060 13.800 1.260 ;
        RECT  12.780 0.800 12.940 1.920 ;
        RECT  11.500 1.760 12.940 1.920 ;
        RECT  11.300 0.300 12.220 0.460 ;
        RECT  12.060 0.300 12.220 0.640 ;
        RECT  12.060 0.480 13.330 0.640 ;
        RECT  13.170 0.480 13.330 0.860 ;
        RECT  13.170 0.700 14.240 0.860 ;
        RECT  10.380 0.580 10.560 1.780 ;
        RECT  11.300 0.300 11.460 1.150 ;
        RECT  10.380 0.990 11.460 1.150 ;
        RECT  14.720 1.060 15.820 1.260 ;
        RECT  13.220 1.420 14.240 1.580 ;
        RECT  10.380 0.990 10.580 1.780 ;
        RECT  14.080 0.700 14.240 2.100 ;
        RECT  13.220 1.420 13.420 2.000 ;
        RECT  14.720 1.060 14.880 2.100 ;
        RECT  14.080 1.940 14.880 2.100 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  8.760 0.900 8.960 1.100 ;
        LAYER ME2 ;
        RECT  6.720 0.400 8.960 0.600 ;
        RECT  8.760 0.400 8.960 1.200 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.090 2.400 ;
        RECT  0.000 1.160 5.660 2.400 ;
        RECT  7.070 1.080 9.930 2.400 ;
        RECT  10.800 1.140 16.400 2.400 ;
        RECT  0.000 1.200 16.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.400 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.930 0.000 16.400 1.140 ;
        RECT  4.090 0.000 7.070 1.160 ;
        RECT  5.660 0.000 7.070 1.200 ;
        RECT  9.930 0.000 10.800 1.200 ;
    END
END SDFSM4HM

MACRO SDFSM2HM
    CLASS CORE ;
    FOREIGN SDFSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.516  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 0.940 2.860 1.340 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.160 0.840 3.500 1.220 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.480 1.460 14.300 1.640 ;
        RECT  14.100 0.740 14.300 1.640 ;
        RECT  13.480 0.740 14.300 0.900 ;
        RECT  13.480 1.460 13.640 1.950 ;
        RECT  13.480 0.400 13.640 0.900 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.420 1.880 14.700 2.080 ;
        RECT  14.500 0.350 14.700 2.080 ;
        RECT  14.420 0.350 14.700 0.550 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.192  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.700 1.430 11.920 1.590 ;
        RECT  11.640 1.120 11.920 1.590 ;
        RECT  10.080 1.940 10.860 2.100 ;
        RECT  10.700 1.430 10.860 2.100 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  13.940 1.840 14.140 2.540 ;
        RECT  12.810 2.080 13.090 2.540 ;
        RECT  11.980 2.080 12.260 2.540 ;
        RECT  11.020 1.840 11.220 2.540 ;
        RECT  7.980 2.080 8.260 2.540 ;
        RECT  4.320 2.020 4.520 2.540 ;
        RECT  2.940 1.980 3.100 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  13.940 -0.140 14.140 0.560 ;
        RECT  12.900 -0.140 13.180 0.500 ;
        RECT  10.940 -0.140 11.100 0.650 ;
        RECT  7.360 -0.140 7.560 0.560 ;
        RECT  4.420 -0.140 4.620 0.600 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.700 ;
        RECT  2.160 1.500 2.460 1.700 ;
        RECT  3.660 0.620 3.940 1.300 ;
        RECT  3.660 1.100 4.780 1.300 ;
        RECT  3.660 0.620 3.820 1.760 ;
        RECT  2.620 1.660 3.420 1.820 ;
        RECT  3.980 1.700 4.840 1.860 ;
        RECT  3.260 1.660 3.420 2.100 ;
        RECT  4.680 1.700 4.840 2.100 ;
        RECT  2.620 1.660 2.780 2.020 ;
        RECT  1.580 1.860 2.780 2.020 ;
        RECT  3.980 1.700 4.160 2.100 ;
        RECT  3.260 1.940 4.160 2.100 ;
        RECT  5.480 1.740 5.680 2.100 ;
        RECT  4.680 1.940 5.680 2.100 ;
        RECT  1.840 0.300 4.260 0.460 ;
        RECT  4.780 0.300 5.820 0.460 ;
        RECT  5.620 0.300 5.820 0.600 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.100 0.300 4.260 0.920 ;
        RECT  4.780 0.300 4.940 0.920 ;
        RECT  4.100 0.760 4.940 0.920 ;
        RECT  5.980 0.300 6.860 0.460 ;
        RECT  6.660 0.300 6.860 0.720 ;
        RECT  5.100 0.640 5.380 0.920 ;
        RECT  5.980 0.300 6.140 0.920 ;
        RECT  5.100 0.760 6.140 0.920 ;
        RECT  5.100 0.640 5.300 1.510 ;
        RECT  5.000 1.350 5.200 1.780 ;
        RECT  6.300 0.900 7.840 1.060 ;
        RECT  7.640 0.900 7.840 1.220 ;
        RECT  6.300 0.620 6.500 1.400 ;
        RECT  6.000 1.240 6.500 1.400 ;
        RECT  6.000 1.240 6.200 2.020 ;
        RECT  8.000 0.350 8.540 0.550 ;
        RECT  6.880 1.240 7.080 1.600 ;
        RECT  8.000 0.350 8.160 1.600 ;
        RECT  6.880 1.440 8.940 1.600 ;
        RECT  8.740 1.440 8.940 1.780 ;
        RECT  9.100 0.980 9.440 1.180 ;
        RECT  6.360 1.760 8.580 1.920 ;
        RECT  8.420 1.760 8.580 2.100 ;
        RECT  6.360 1.760 6.640 2.100 ;
        RECT  9.100 0.980 9.260 2.100 ;
        RECT  8.420 1.940 9.260 2.100 ;
        RECT  8.720 0.660 9.860 0.820 ;
        RECT  8.720 0.660 8.920 1.200 ;
        RECT  9.700 0.660 9.860 1.270 ;
        RECT  8.820 0.300 10.180 0.500 ;
        RECT  10.020 0.300 10.180 1.760 ;
        RECT  9.420 1.480 10.180 1.760 ;
        RECT  11.580 0.620 11.860 0.960 ;
        RECT  11.580 0.800 12.240 0.960 ;
        RECT  12.080 1.060 13.000 1.260 ;
        RECT  12.080 0.800 12.240 1.920 ;
        RECT  11.460 1.760 12.240 1.920 ;
        RECT  11.260 0.300 12.660 0.460 ;
        RECT  12.100 0.300 12.660 0.590 ;
        RECT  12.500 0.300 12.660 0.900 ;
        RECT  12.500 0.740 13.320 0.900 ;
        RECT  10.340 0.580 10.520 1.780 ;
        RECT  11.260 0.300 11.420 1.150 ;
        RECT  10.340 0.990 11.420 1.150 ;
        RECT  13.160 1.060 13.940 1.260 ;
        RECT  13.160 0.740 13.320 1.580 ;
        RECT  12.460 1.420 13.320 1.580 ;
        RECT  12.460 1.420 12.660 1.720 ;
        RECT  10.340 0.990 10.540 1.780 ;
        LAYER VI1 ;
        RECT  6.660 0.400 6.860 0.600 ;
        RECT  8.720 0.900 8.920 1.100 ;
        LAYER ME2 ;
        RECT  6.560 0.400 8.920 0.600 ;
        RECT  8.720 0.400 8.920 1.200 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.990 2.400 ;
        RECT  0.000 1.160 5.620 2.400 ;
        RECT  6.910 1.080 9.890 2.400 ;
        RECT  10.760 1.140 14.800 2.400 ;
        RECT  0.000 1.200 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.080 ;
        RECT  0.000 0.000 6.910 1.140 ;
        RECT  9.890 0.000 14.800 1.140 ;
        RECT  3.990 0.000 6.910 1.160 ;
        RECT  5.620 0.000 6.910 1.200 ;
        RECT  9.890 0.000 10.760 1.200 ;
    END
END SDFSM2HM

MACRO SDFSM1HM
    CLASS CORE ;
    FOREIGN SDFSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.344  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.000 0.980 2.200 1.180 ;
        LAYER ME2 ;
        RECT  2.000 0.820 2.300 1.330 ;
        LAYER ME1 ;
        RECT  1.920 0.850 2.200 1.280 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.840 3.190 1.300 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.400 1.460 14.300 1.660 ;
        RECT  14.100 0.740 14.300 1.660 ;
        RECT  13.400 0.740 14.300 0.900 ;
        RECT  13.400 1.460 13.600 2.000 ;
        RECT  13.400 0.350 13.600 0.900 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.360 1.850 14.700 2.050 ;
        RECT  14.500 0.350 14.700 2.050 ;
        RECT  14.360 0.350 14.700 0.550 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.172  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.560 1.430 11.900 1.590 ;
        RECT  11.620 1.120 11.900 1.590 ;
        RECT  9.940 1.940 10.720 2.100 ;
        RECT  10.560 1.430 10.720 2.100 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  13.880 1.840 14.080 2.540 ;
        RECT  12.820 2.020 13.020 2.540 ;
        RECT  11.840 2.080 12.120 2.540 ;
        RECT  10.880 1.840 11.080 2.540 ;
        RECT  7.840 2.080 8.120 2.540 ;
        RECT  4.180 1.780 4.380 2.540 ;
        RECT  2.640 2.080 2.920 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  13.880 -0.140 14.080 0.560 ;
        RECT  12.840 -0.140 13.120 0.500 ;
        RECT  10.800 -0.140 10.960 0.650 ;
        RECT  7.220 -0.140 7.420 0.560 ;
        RECT  4.180 -0.140 4.380 0.600 ;
        RECT  2.660 -0.140 2.940 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.440 2.680 1.600 ;
        RECT  2.480 0.850 2.680 1.600 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  3.420 0.620 3.700 0.840 ;
        RECT  3.540 1.080 4.640 1.280 ;
        RECT  3.540 0.620 3.700 1.780 ;
        RECT  3.860 1.460 4.700 1.620 ;
        RECT  1.950 1.760 3.240 1.920 ;
        RECT  3.080 1.760 3.240 2.100 ;
        RECT  4.540 1.460 4.700 2.100 ;
        RECT  1.580 1.860 2.100 2.020 ;
        RECT  3.860 1.460 4.020 2.100 ;
        RECT  3.080 1.940 4.020 2.100 ;
        RECT  5.340 1.740 5.540 2.100 ;
        RECT  4.540 1.940 5.540 2.100 ;
        RECT  3.100 0.300 4.020 0.460 ;
        RECT  4.540 0.300 5.580 0.460 ;
        RECT  1.820 0.360 2.020 0.640 ;
        RECT  5.380 0.300 5.580 0.600 ;
        RECT  3.100 0.300 3.260 0.640 ;
        RECT  1.820 0.480 3.260 0.640 ;
        RECT  3.860 0.300 4.020 0.920 ;
        RECT  4.540 0.300 4.700 0.920 ;
        RECT  3.860 0.760 4.700 0.920 ;
        RECT  5.740 0.300 6.620 0.460 ;
        RECT  6.420 0.300 6.620 0.720 ;
        RECT  4.860 0.620 5.140 0.920 ;
        RECT  5.740 0.300 5.900 0.920 ;
        RECT  4.860 0.760 5.900 0.920 ;
        RECT  4.860 0.620 5.060 1.780 ;
        RECT  6.060 0.900 7.700 1.060 ;
        RECT  7.500 0.900 7.700 1.220 ;
        RECT  6.060 0.620 6.260 1.400 ;
        RECT  5.860 1.240 6.060 2.020 ;
        RECT  7.860 0.350 8.400 0.550 ;
        RECT  6.740 1.240 6.940 1.600 ;
        RECT  7.860 0.350 8.020 1.600 ;
        RECT  6.740 1.440 8.800 1.600 ;
        RECT  8.600 1.440 8.800 1.780 ;
        RECT  8.960 0.980 9.300 1.180 ;
        RECT  6.220 1.760 8.440 1.920 ;
        RECT  8.280 1.760 8.440 2.100 ;
        RECT  6.220 1.760 6.500 2.100 ;
        RECT  8.960 0.980 9.120 2.100 ;
        RECT  8.280 1.940 9.120 2.100 ;
        RECT  8.580 0.660 9.720 0.820 ;
        RECT  8.580 0.660 8.780 1.200 ;
        RECT  9.560 0.660 9.720 1.270 ;
        RECT  8.680 0.300 10.040 0.500 ;
        RECT  9.880 0.300 10.040 1.760 ;
        RECT  9.280 1.480 10.040 1.760 ;
        RECT  11.440 0.620 11.720 0.960 ;
        RECT  11.440 0.800 12.220 0.960 ;
        RECT  12.060 1.060 12.900 1.260 ;
        RECT  12.060 0.800 12.220 1.920 ;
        RECT  11.320 1.760 12.220 1.920 ;
        RECT  11.120 0.300 12.580 0.460 ;
        RECT  11.960 0.300 12.580 0.580 ;
        RECT  12.420 0.300 12.580 0.900 ;
        RECT  12.420 0.740 13.220 0.900 ;
        RECT  10.200 0.580 10.380 1.780 ;
        RECT  11.120 0.300 11.280 1.150 ;
        RECT  10.200 0.990 11.280 1.150 ;
        RECT  13.060 1.060 13.900 1.260 ;
        RECT  13.060 0.740 13.220 1.580 ;
        RECT  12.380 1.420 13.220 1.580 ;
        RECT  10.200 0.990 10.400 1.780 ;
        RECT  12.380 1.420 12.540 1.780 ;
        LAYER VI1 ;
        RECT  6.420 0.400 6.620 0.600 ;
        RECT  8.580 0.900 8.780 1.100 ;
        LAYER ME2 ;
        RECT  6.320 0.400 8.780 0.600 ;
        RECT  8.580 0.400 8.780 1.200 ;
        LAYER VTPH ;
        RECT  1.540 1.050 2.670 2.400 ;
        RECT  0.000 1.140 2.670 2.400 ;
        RECT  0.000 1.160 5.480 2.400 ;
        RECT  6.670 1.080 9.750 2.400 ;
        RECT  10.600 1.140 14.800 2.400 ;
        RECT  0.000 1.200 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.050 ;
        RECT  2.670 0.000 14.800 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  9.750 0.000 14.800 1.140 ;
        RECT  2.670 0.000 6.670 1.160 ;
        RECT  5.480 0.000 6.670 1.200 ;
        RECT  9.750 0.000 10.600 1.200 ;
    END
END SDFSM1HM

MACRO SDFRSM8HM
    CLASS CORE ;
    FOREIGN SDFRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.190 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.314  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.700 0.410 17.860 1.780 ;
        RECT  16.420 0.850 17.860 1.100 ;
        RECT  16.420 0.410 16.580 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  19.880 0.450 20.080 2.080 ;
        RECT  18.840 1.440 20.080 1.630 ;
        RECT  19.700 0.660 20.080 1.630 ;
        RECT  18.840 0.660 20.080 0.820 ;
        RECT  18.840 1.440 19.040 2.080 ;
        RECT  18.840 0.450 19.040 0.820 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.319  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 9.810  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.980 0.800 13.260 1.060 ;
        RECT  12.000 0.800 13.260 0.960 ;
        RECT  12.000 0.800 12.300 1.240 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.234  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.990 0.900 15.560 1.160 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 20.800 2.540 ;
        RECT  20.400 1.480 20.600 2.540 ;
        RECT  19.320 1.900 19.600 2.540 ;
        RECT  18.340 1.440 18.500 2.540 ;
        RECT  17.060 1.800 17.220 2.540 ;
        RECT  15.740 2.020 15.940 2.540 ;
        RECT  14.540 1.860 14.820 2.540 ;
        RECT  13.400 1.860 13.680 2.540 ;
        RECT  12.320 1.800 12.520 2.540 ;
        RECT  8.920 2.080 9.200 2.540 ;
        RECT  4.360 1.980 4.520 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 20.800 0.140 ;
        RECT  20.400 -0.140 20.600 0.730 ;
        RECT  19.320 -0.140 19.600 0.500 ;
        RECT  18.320 -0.140 18.520 0.730 ;
        RECT  17.040 -0.140 17.240 0.560 ;
        RECT  15.700 -0.140 15.980 0.320 ;
        RECT  14.340 -0.140 14.620 0.320 ;
        RECT  12.220 -0.140 12.500 0.320 ;
        RECT  7.900 -0.140 8.100 0.400 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.300 ;
        RECT  3.700 1.100 4.820 1.300 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.660 4.840 1.820 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.680 1.660 4.840 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.660 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.680 1.940 5.660 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.640 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.640 5.460 1.510 ;
        RECT  5.000 1.350 5.460 1.510 ;
        RECT  5.000 1.350 5.160 1.780 ;
        RECT  6.720 1.620 8.160 1.780 ;
        RECT  6.460 0.900 8.800 1.060 ;
        RECT  8.640 0.900 8.800 1.260 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  5.980 1.240 6.660 1.400 ;
        RECT  5.980 1.240 6.180 2.020 ;
        RECT  8.960 0.620 9.700 0.780 ;
        RECT  6.930 1.240 8.480 1.400 ;
        RECT  8.320 1.240 8.480 1.600 ;
        RECT  8.960 0.620 9.120 1.600 ;
        RECT  8.320 1.440 9.880 1.600 ;
        RECT  9.680 1.440 9.880 1.760 ;
        RECT  8.320 1.760 9.520 1.920 ;
        RECT  9.360 1.760 9.520 2.100 ;
        RECT  8.320 1.760 8.480 2.100 ;
        RECT  6.340 1.940 8.480 2.100 ;
        RECT  10.080 1.660 10.240 2.100 ;
        RECT  9.360 1.940 10.240 2.100 ;
        RECT  9.720 1.080 11.200 1.280 ;
        RECT  8.260 0.300 11.240 0.460 ;
        RECT  7.460 0.300 7.740 0.720 ;
        RECT  8.260 0.300 8.420 0.720 ;
        RECT  7.460 0.560 8.420 0.720 ;
        RECT  10.020 0.620 10.300 0.900 ;
        RECT  10.020 0.740 11.520 0.900 ;
        RECT  12.460 1.120 12.780 1.380 ;
        RECT  14.120 1.120 14.400 1.380 ;
        RECT  12.460 1.220 14.400 1.380 ;
        RECT  12.460 1.120 12.620 1.640 ;
        RECT  12.000 1.480 12.620 1.640 ;
        RECT  10.780 1.510 11.520 1.710 ;
        RECT  11.360 0.740 11.520 2.100 ;
        RECT  11.350 1.510 11.520 2.100 ;
        RECT  12.000 1.480 12.160 2.100 ;
        RECT  11.350 1.940 12.160 2.100 ;
        RECT  13.420 0.620 13.700 0.960 ;
        RECT  13.420 0.800 14.720 0.960 ;
        RECT  15.780 0.980 15.940 1.480 ;
        RECT  14.560 1.320 15.940 1.480 ;
        RECT  14.560 0.800 14.720 1.700 ;
        RECT  12.800 1.540 14.720 1.700 ;
        RECT  12.660 0.300 14.100 0.460 ;
        RECT  13.940 0.300 14.100 0.640 ;
        RECT  12.660 0.300 12.820 0.640 ;
        RECT  11.680 0.480 12.820 0.640 ;
        RECT  13.940 0.480 16.260 0.640 ;
        RECT  18.020 1.020 19.260 1.220 ;
        RECT  16.740 1.480 17.540 1.640 ;
        RECT  11.680 0.480 11.840 1.780 ;
        RECT  15.020 1.700 16.260 1.860 ;
        RECT  16.100 0.480 16.260 2.100 ;
        RECT  17.380 1.480 17.540 2.100 ;
        RECT  16.740 1.480 16.900 2.100 ;
        RECT  16.100 1.940 16.900 2.100 ;
        RECT  18.020 1.020 18.180 2.100 ;
        RECT  17.380 1.940 18.180 2.100 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  9.820 1.080 10.020 1.280 ;
        LAYER ME2 ;
        RECT  6.720 0.400 10.020 0.600 ;
        RECT  9.820 0.400 10.020 1.380 ;
        LAYER VTPH ;
        RECT  7.070 1.080 9.200 2.400 ;
        RECT  12.220 1.080 13.070 2.400 ;
        RECT  0.000 1.140 4.090 2.400 ;
        RECT  0.000 1.160 5.660 2.400 ;
        RECT  7.070 1.140 20.800 2.400 ;
        RECT  0.000 1.200 20.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 20.800 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.200 0.000 12.220 1.140 ;
        RECT  13.070 0.000 20.800 1.140 ;
        RECT  4.090 0.000 7.070 1.160 ;
        RECT  5.660 0.000 7.070 1.200 ;
    END
END SDFRSM8HM

MACRO SDFRSM4HM
    CLASS CORE ;
    FOREIGN SDFRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.319  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 16.953  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 19.538  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  12.020 0.760 12.220 0.960 ;
        LAYER ME2 ;
        RECT  12.020 0.660 12.300 1.160 ;
        LAYER ME1 ;
        RECT  12.000 0.620 12.240 1.060 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.670  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.400 0.850 15.960 1.150 ;
        RECT  15.400 0.410 15.560 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.540 1.440 17.100 1.640 ;
        RECT  16.900 0.660 17.100 1.640 ;
        RECT  16.540 0.660 17.100 0.820 ;
        RECT  16.540 1.440 16.740 2.080 ;
        RECT  16.540 0.450 16.740 0.820 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.241  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.970 0.900 14.390 1.160 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.600 2.540 ;
        RECT  17.060 1.840 17.260 2.540 ;
        RECT  16.040 1.800 16.200 2.540 ;
        RECT  14.720 2.020 14.920 2.540 ;
        RECT  13.520 1.860 13.800 2.540 ;
        RECT  12.380 1.580 12.660 2.540 ;
        RECT  8.920 2.080 9.200 2.540 ;
        RECT  4.360 1.980 4.520 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.600 0.140 ;
        RECT  17.020 -0.140 17.300 0.500 ;
        RECT  16.020 -0.140 16.220 0.560 ;
        RECT  14.680 -0.140 14.960 0.320 ;
        RECT  13.320 -0.140 13.600 0.320 ;
        RECT  7.900 -0.140 8.100 0.400 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.300 ;
        RECT  3.700 1.100 4.820 1.300 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.660 4.840 1.820 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.680 1.660 4.840 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.660 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.680 1.940 5.660 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.640 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.640 5.460 1.510 ;
        RECT  5.000 1.350 5.460 1.510 ;
        RECT  5.000 1.350 5.160 1.780 ;
        RECT  6.720 1.620 8.160 1.780 ;
        RECT  6.460 0.900 8.800 1.060 ;
        RECT  8.640 0.900 8.800 1.260 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  5.980 1.240 6.660 1.400 ;
        RECT  5.980 1.240 6.180 2.020 ;
        RECT  8.960 0.620 9.700 0.780 ;
        RECT  6.930 1.240 8.480 1.400 ;
        RECT  8.320 1.240 8.480 1.600 ;
        RECT  8.960 0.620 9.120 1.600 ;
        RECT  8.320 1.440 9.880 1.600 ;
        RECT  9.680 1.440 9.880 1.760 ;
        RECT  8.320 1.760 9.520 1.920 ;
        RECT  9.360 1.760 9.520 2.100 ;
        RECT  8.320 1.760 8.480 2.100 ;
        RECT  6.340 1.940 8.480 2.100 ;
        RECT  10.080 1.660 10.240 2.100 ;
        RECT  9.360 1.940 10.240 2.100 ;
        RECT  9.720 1.080 11.200 1.280 ;
        RECT  8.260 0.300 11.240 0.460 ;
        RECT  7.460 0.300 7.740 0.720 ;
        RECT  8.260 0.300 8.420 0.720 ;
        RECT  7.460 0.560 8.420 0.720 ;
        RECT  10.020 0.620 10.300 0.900 ;
        RECT  10.020 0.740 11.520 0.900 ;
        RECT  13.100 1.120 13.380 1.380 ;
        RECT  12.000 1.220 13.380 1.380 ;
        RECT  10.780 1.510 11.520 1.710 ;
        RECT  11.360 0.740 11.520 2.100 ;
        RECT  11.350 1.510 11.520 2.100 ;
        RECT  12.000 1.220 12.160 2.100 ;
        RECT  11.350 1.940 12.160 2.100 ;
        RECT  12.400 0.620 12.680 0.960 ;
        RECT  12.400 0.800 13.700 0.960 ;
        RECT  14.760 0.980 14.920 1.480 ;
        RECT  13.540 1.320 14.920 1.480 ;
        RECT  13.540 0.800 13.700 1.700 ;
        RECT  12.920 1.540 13.700 1.700 ;
        RECT  11.680 0.300 13.080 0.460 ;
        RECT  12.920 0.300 13.080 0.640 ;
        RECT  12.920 0.480 15.240 0.640 ;
        RECT  16.120 1.020 16.600 1.220 ;
        RECT  16.120 1.020 16.280 1.640 ;
        RECT  15.720 1.480 16.280 1.640 ;
        RECT  11.680 0.300 11.840 1.780 ;
        RECT  14.000 1.700 15.240 1.860 ;
        RECT  15.080 0.480 15.240 2.100 ;
        RECT  15.720 1.480 15.880 2.100 ;
        RECT  15.080 1.940 15.880 2.100 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  9.820 1.080 10.020 1.280 ;
        LAYER ME2 ;
        RECT  6.720 0.400 10.020 0.600 ;
        RECT  9.820 0.400 10.020 1.380 ;
        LAYER VTPH ;
        RECT  7.070 1.080 9.200 2.400 ;
        RECT  0.000 1.140 4.090 2.400 ;
        RECT  0.000 1.160 5.660 2.400 ;
        RECT  7.070 1.140 17.600 2.400 ;
        RECT  0.000 1.200 17.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.600 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.200 0.000 17.600 1.140 ;
        RECT  4.090 0.000 7.070 1.160 ;
        RECT  5.660 0.000 7.070 1.200 ;
    END
END SDFRSM4HM

MACRO SDFRSM2HM
    CLASS CORE ;
    FOREIGN SDFRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.184  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.970 0.830 14.390 1.100 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.319  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 16.953  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 19.538  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  12.020 0.760 12.220 0.960 ;
        LAYER ME2 ;
        RECT  12.020 0.660 12.300 1.160 ;
        LAYER ME1 ;
        RECT  12.000 0.620 12.240 1.060 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.583  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.400 1.460 16.300 1.660 ;
        RECT  16.100 0.670 16.300 1.660 ;
        RECT  15.410 0.670 16.300 0.830 ;
        RECT  15.400 1.460 15.610 2.100 ;
        RECT  15.410 0.380 15.610 0.830 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.460 0.450 16.700 2.080 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.800 2.540 ;
        RECT  15.940 1.840 16.140 2.540 ;
        RECT  14.720 2.020 14.920 2.540 ;
        RECT  13.520 1.860 13.800 2.540 ;
        RECT  12.380 1.580 12.660 2.540 ;
        RECT  8.920 2.080 9.200 2.540 ;
        RECT  4.360 1.980 4.520 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.800 0.140 ;
        RECT  15.900 -0.140 16.180 0.500 ;
        RECT  14.680 -0.140 14.960 0.320 ;
        RECT  13.320 -0.140 13.600 0.320 ;
        RECT  7.900 -0.140 8.100 0.400 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.300 ;
        RECT  3.700 1.100 4.820 1.300 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.660 4.840 1.820 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.680 1.660 4.840 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.660 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.680 1.940 5.660 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.640 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.640 5.460 1.510 ;
        RECT  5.000 1.350 5.460 1.510 ;
        RECT  5.000 1.350 5.160 1.780 ;
        RECT  6.720 1.620 8.160 1.780 ;
        RECT  6.460 0.900 8.800 1.060 ;
        RECT  8.640 0.900 8.800 1.260 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  5.980 1.240 6.660 1.400 ;
        RECT  5.980 1.240 6.180 2.020 ;
        RECT  8.960 0.620 9.700 0.780 ;
        RECT  6.930 1.240 8.480 1.400 ;
        RECT  8.320 1.240 8.480 1.600 ;
        RECT  8.960 0.620 9.120 1.600 ;
        RECT  8.320 1.440 9.880 1.600 ;
        RECT  9.680 1.440 9.880 1.760 ;
        RECT  8.320 1.760 9.520 1.920 ;
        RECT  9.360 1.760 9.520 2.100 ;
        RECT  8.320 1.760 8.480 2.100 ;
        RECT  6.340 1.940 8.480 2.100 ;
        RECT  10.080 1.660 10.240 2.100 ;
        RECT  9.360 1.940 10.240 2.100 ;
        RECT  9.720 1.080 11.200 1.280 ;
        RECT  8.260 0.300 11.240 0.460 ;
        RECT  7.460 0.300 7.740 0.720 ;
        RECT  8.260 0.300 8.420 0.720 ;
        RECT  7.460 0.560 8.420 0.720 ;
        RECT  10.020 0.620 10.300 0.900 ;
        RECT  10.020 0.740 11.520 0.900 ;
        RECT  13.100 1.120 13.380 1.380 ;
        RECT  12.000 1.220 13.380 1.380 ;
        RECT  10.780 1.510 11.520 1.710 ;
        RECT  11.360 0.740 11.520 2.100 ;
        RECT  11.350 1.510 11.520 2.100 ;
        RECT  12.000 1.220 12.160 2.100 ;
        RECT  11.350 1.940 12.160 2.100 ;
        RECT  12.400 0.620 12.680 0.960 ;
        RECT  12.400 0.800 13.700 0.960 ;
        RECT  14.550 1.060 14.750 1.420 ;
        RECT  13.540 1.260 14.750 1.420 ;
        RECT  13.540 0.800 13.700 1.700 ;
        RECT  12.920 1.540 13.700 1.700 ;
        RECT  11.680 0.300 13.080 0.460 ;
        RECT  12.920 0.300 13.080 0.640 ;
        RECT  12.920 0.480 15.240 0.640 ;
        RECT  15.080 1.020 15.880 1.220 ;
        RECT  11.680 0.300 11.840 1.780 ;
        RECT  15.080 0.480 15.240 1.860 ;
        RECT  14.040 1.700 15.240 1.860 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  9.820 1.080 10.020 1.280 ;
        LAYER ME2 ;
        RECT  6.720 0.400 10.020 0.600 ;
        RECT  9.820 0.400 10.020 1.380 ;
        LAYER VTPH ;
        RECT  7.070 1.080 9.200 2.400 ;
        RECT  0.000 1.140 4.090 2.400 ;
        RECT  0.000 1.160 5.660 2.400 ;
        RECT  7.070 1.140 16.800 2.400 ;
        RECT  0.000 1.200 16.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.800 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.200 0.000 16.800 1.140 ;
        RECT  4.090 0.000 7.070 1.160 ;
        RECT  5.660 0.000 7.070 1.200 ;
    END
END SDFRSM2HM

MACRO SDFRSM1HM
    CLASS CORE ;
    FOREIGN SDFRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.344  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.930 0.960 2.130 1.160 ;
        LAYER ME2 ;
        RECT  1.930 0.840 2.300 1.280 ;
        LAYER ME1 ;
        RECT  1.800 0.900 2.190 1.220 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.840 3.160 1.300 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.343  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.120 0.440 15.500 0.760 ;
        RECT  15.120 0.440 15.280 1.760 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.100 1.570 16.500 1.770 ;
        RECT  16.100 0.420 16.500 0.620 ;
        RECT  16.100 0.420 16.300 1.770 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.345  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 17.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.720 0.800 12.880 1.240 ;
        RECT  11.700 0.800 12.880 0.960 ;
        RECT  11.700 0.800 11.980 1.160 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.640 1.160 13.960 1.500 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.870 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.800 2.540 ;
        RECT  15.760 1.490 15.920 2.540 ;
        RECT  14.300 2.020 14.500 2.540 ;
        RECT  13.080 1.860 13.360 2.540 ;
        RECT  12.000 1.800 12.200 2.540 ;
        RECT  8.550 2.080 8.830 2.540 ;
        RECT  4.150 2.020 4.350 2.540 ;
        RECT  2.680 2.020 2.880 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.800 0.140 ;
        RECT  15.740 -0.140 15.940 0.660 ;
        RECT  14.500 -0.140 14.780 0.320 ;
        RECT  11.890 -0.140 12.170 0.320 ;
        RECT  7.530 -0.140 7.810 0.420 ;
        RECT  4.130 -0.140 4.330 0.600 ;
        RECT  2.660 -0.140 2.940 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.380 2.680 1.540 ;
        RECT  2.480 0.850 2.680 1.540 ;
        RECT  1.440 1.070 1.640 1.700 ;
        RECT  0.140 1.540 1.640 1.700 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  3.420 1.100 4.610 1.300 ;
        RECT  3.420 0.620 3.620 1.780 ;
        RECT  1.950 1.700 3.200 1.860 ;
        RECT  3.810 1.700 4.670 1.860 ;
        RECT  3.040 1.700 3.200 2.100 ;
        RECT  4.510 1.700 4.670 2.100 ;
        RECT  1.580 1.860 2.110 2.020 ;
        RECT  3.810 1.700 3.990 2.100 ;
        RECT  3.040 1.940 3.990 2.100 ;
        RECT  5.310 1.740 5.510 2.100 ;
        RECT  4.510 1.940 5.510 2.100 ;
        RECT  3.100 0.300 3.970 0.460 ;
        RECT  4.490 0.300 5.550 0.460 ;
        RECT  1.820 0.370 2.020 0.680 ;
        RECT  5.350 0.300 5.550 0.600 ;
        RECT  3.100 0.300 3.260 0.680 ;
        RECT  1.820 0.520 3.260 0.680 ;
        RECT  3.810 0.300 3.970 0.920 ;
        RECT  4.490 0.300 4.650 0.920 ;
        RECT  3.810 0.760 4.650 0.920 ;
        RECT  5.710 0.300 6.670 0.460 ;
        RECT  6.470 0.300 6.670 0.720 ;
        RECT  4.830 0.640 5.110 0.920 ;
        RECT  5.710 0.300 5.870 0.920 ;
        RECT  4.830 0.760 5.870 0.920 ;
        RECT  4.830 0.640 5.030 1.780 ;
        RECT  6.390 1.560 7.750 1.780 ;
        RECT  6.030 0.920 7.950 1.080 ;
        RECT  6.030 0.680 6.310 1.400 ;
        RECT  5.830 1.240 6.030 2.020 ;
        RECT  8.630 0.620 9.330 0.780 ;
        RECT  6.710 1.240 8.110 1.400 ;
        RECT  7.950 1.240 8.110 1.600 ;
        RECT  8.630 0.620 8.790 1.600 ;
        RECT  7.950 1.440 9.520 1.600 ;
        RECT  9.320 1.440 9.520 1.780 ;
        RECT  7.950 1.760 9.160 1.920 ;
        RECT  9.000 1.760 9.160 2.100 ;
        RECT  7.950 1.760 8.110 2.100 ;
        RECT  6.190 1.940 8.110 2.100 ;
        RECT  9.720 1.660 9.880 2.100 ;
        RECT  9.000 1.940 9.880 2.100 ;
        RECT  9.350 1.080 10.840 1.280 ;
        RECT  7.970 0.300 10.880 0.460 ;
        RECT  7.090 0.300 7.370 0.740 ;
        RECT  7.970 0.300 8.130 0.740 ;
        RECT  7.090 0.580 8.130 0.740 ;
        RECT  9.710 0.620 9.990 0.900 ;
        RECT  9.710 0.740 11.160 0.900 ;
        RECT  12.180 1.120 12.460 1.340 ;
        RECT  11.680 1.320 12.340 1.480 ;
        RECT  10.460 1.460 10.660 1.920 ;
        RECT  10.460 1.760 11.160 1.920 ;
        RECT  11.000 0.740 11.160 2.100 ;
        RECT  10.990 1.760 11.160 2.100 ;
        RECT  11.680 1.320 11.840 2.100 ;
        RECT  10.990 1.940 11.840 2.100 ;
        RECT  13.040 0.620 13.360 0.960 ;
        RECT  13.040 0.800 14.500 0.960 ;
        RECT  14.300 0.800 14.500 1.300 ;
        RECT  13.040 0.620 13.200 1.700 ;
        RECT  12.520 1.500 13.200 1.700 ;
        RECT  12.330 0.300 13.800 0.460 ;
        RECT  13.600 0.300 13.800 0.640 ;
        RECT  12.330 0.300 12.490 0.640 ;
        RECT  11.320 0.480 12.490 0.640 ;
        RECT  13.600 0.480 14.820 0.640 ;
        RECT  15.440 1.020 15.880 1.220 ;
        RECT  11.320 0.480 11.520 1.760 ;
        RECT  13.640 1.700 14.820 1.860 ;
        RECT  14.660 0.480 14.820 2.100 ;
        RECT  15.440 1.020 15.600 2.100 ;
        RECT  14.660 1.940 15.600 2.100 ;
        LAYER VI1 ;
        RECT  6.470 0.400 6.670 0.600 ;
        RECT  9.450 1.080 9.650 1.280 ;
        LAYER ME2 ;
        RECT  6.370 0.400 9.650 0.600 ;
        RECT  9.450 0.400 9.650 1.380 ;
        LAYER VTPH ;
        RECT  7.480 1.080 8.830 2.400 ;
        RECT  1.370 1.050 2.650 2.400 ;
        RECT  0.000 1.140 2.650 2.400 ;
        RECT  7.480 1.140 16.800 2.400 ;
        RECT  0.000 1.200 16.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.800 1.050 ;
        RECT  2.650 0.000 16.800 1.080 ;
        RECT  0.000 0.000 1.370 1.140 ;
        RECT  8.830 0.000 16.800 1.140 ;
        RECT  2.650 0.000 7.480 1.200 ;
    END
END SDFRSM1HM

MACRO SDFRM8HM
    CLASS CORE ;
    FOREIGN SDFRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.481  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.010 2.860 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.190 1.050 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.166  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.200 1.440 16.800 1.600 ;
        RECT  15.320 0.660 16.720 0.820 ;
        RECT  16.520 0.430 16.720 0.820 ;
        RECT  16.100 0.660 16.300 1.600 ;
        RECT  15.320 0.430 15.520 0.820 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  18.720 1.440 19.030 2.080 ;
        RECT  17.680 0.660 19.030 0.860 ;
        RECT  18.720 0.430 19.030 0.860 ;
        RECT  17.680 1.440 19.030 1.640 ;
        RECT  18.500 0.660 18.700 1.640 ;
        RECT  17.680 1.440 17.880 2.080 ;
        RECT  17.680 0.430 17.880 0.860 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.830 1.120 13.490 1.280 ;
        RECT  11.830 0.900 12.360 1.280 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 19.600 2.540 ;
        RECT  19.240 1.480 19.440 2.540 ;
        RECT  18.200 1.840 18.400 2.540 ;
        RECT  17.080 2.080 17.360 2.540 ;
        RECT  15.880 2.080 16.160 2.540 ;
        RECT  14.670 2.080 14.950 2.540 ;
        RECT  13.590 1.840 13.790 2.540 ;
        RECT  12.510 1.760 12.790 2.540 ;
        RECT  11.730 1.500 11.890 2.540 ;
        RECT  11.450 1.500 11.890 1.700 ;
        RECT  8.700 2.080 8.980 2.540 ;
        RECT  4.360 2.020 4.560 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 19.600 0.140 ;
        RECT  19.240 -0.140 19.440 0.710 ;
        RECT  18.160 -0.140 18.440 0.500 ;
        RECT  17.160 -0.140 17.360 0.710 ;
        RECT  15.880 -0.140 16.160 0.500 ;
        RECT  14.710 -0.140 14.910 0.560 ;
        RECT  13.510 -0.140 13.790 0.320 ;
        RECT  11.070 -0.140 11.350 0.540 ;
        RECT  8.070 -0.140 8.350 0.710 ;
        RECT  4.660 -0.140 4.860 0.610 ;
        RECT  3.140 -0.140 3.420 0.500 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.700 ;
        RECT  0.140 1.540 1.640 1.700 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.900 0.620 4.180 1.300 ;
        RECT  3.720 1.100 4.770 1.300 ;
        RECT  3.720 1.100 3.880 1.760 ;
        RECT  4.040 1.700 4.880 1.860 ;
        RECT  2.600 1.760 3.520 1.920 ;
        RECT  1.620 1.860 1.910 2.100 ;
        RECT  3.360 1.760 3.520 2.100 ;
        RECT  4.720 1.700 4.880 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.040 1.700 4.200 2.100 ;
        RECT  3.360 1.940 4.200 2.100 ;
        RECT  5.520 1.740 5.720 2.100 ;
        RECT  4.720 1.940 5.720 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.580 0.300 4.500 0.460 ;
        RECT  5.020 0.300 6.060 0.460 ;
        RECT  5.860 0.300 6.060 0.600 ;
        RECT  2.820 0.300 2.980 0.820 ;
        RECT  1.840 0.300 2.000 0.690 ;
        RECT  4.340 0.300 4.500 0.930 ;
        RECT  3.580 0.300 3.740 0.820 ;
        RECT  2.820 0.660 3.740 0.820 ;
        RECT  5.020 0.300 5.180 0.930 ;
        RECT  4.340 0.770 5.180 0.930 ;
        RECT  6.220 0.300 7.100 0.460 ;
        RECT  6.900 0.300 7.100 0.700 ;
        RECT  5.340 0.660 5.620 0.920 ;
        RECT  6.220 0.300 6.380 0.920 ;
        RECT  5.340 0.760 6.380 0.920 ;
        RECT  5.340 0.660 5.540 1.450 ;
        RECT  5.040 1.250 5.540 1.450 ;
        RECT  5.040 1.250 5.240 1.780 ;
        RECT  6.780 1.620 8.220 1.780 ;
        RECT  6.540 0.980 8.320 1.140 ;
        RECT  6.540 0.620 6.740 1.240 ;
        RECT  6.040 1.080 6.740 1.240 ;
        RECT  6.040 1.080 6.240 2.020 ;
        RECT  8.800 0.600 9.000 1.600 ;
        RECT  7.160 1.300 9.000 1.460 ;
        RECT  8.800 1.440 9.660 1.600 ;
        RECT  9.460 1.440 9.660 1.780 ;
        RECT  8.380 1.760 9.300 1.920 ;
        RECT  9.140 1.760 9.300 2.100 ;
        RECT  8.380 1.760 8.540 2.100 ;
        RECT  6.400 1.940 8.540 2.100 ;
        RECT  9.140 1.940 9.820 2.100 ;
        RECT  9.440 0.300 10.340 0.460 ;
        RECT  10.180 0.300 10.340 1.310 ;
        RECT  9.440 0.300 9.640 1.280 ;
        RECT  10.180 1.110 10.760 1.310 ;
        RECT  9.820 0.620 10.020 1.780 ;
        RECT  9.820 1.620 10.660 1.780 ;
        RECT  10.490 1.620 10.660 2.100 ;
        RECT  10.490 1.940 11.570 2.100 ;
        RECT  12.470 0.620 12.860 0.780 ;
        RECT  12.700 0.620 12.860 0.960 ;
        RECT  12.700 0.800 14.170 0.960 ;
        RECT  13.970 0.800 14.170 1.600 ;
        RECT  12.050 1.440 14.170 1.600 ;
        RECT  12.050 1.440 12.210 1.840 ;
        RECT  13.070 1.440 13.270 1.870 ;
        RECT  11.510 0.300 13.240 0.460 ;
        RECT  13.080 0.300 13.240 0.640 ;
        RECT  13.080 0.480 14.530 0.640 ;
        RECT  10.500 0.480 10.700 0.860 ;
        RECT  11.510 0.300 11.670 0.860 ;
        RECT  10.500 0.700 11.670 0.860 ;
        RECT  17.050 1.040 18.100 1.240 ;
        RECT  14.370 0.480 14.530 1.920 ;
        RECT  10.980 0.700 11.180 1.780 ;
        RECT  17.050 1.040 17.250 1.920 ;
        RECT  14.070 1.760 17.250 1.920 ;
        LAYER VI1 ;
        RECT  6.900 0.380 7.100 0.580 ;
        RECT  9.440 0.850 9.640 1.050 ;
        LAYER ME2 ;
        RECT  6.750 0.380 9.640 0.580 ;
        RECT  9.440 0.380 9.640 1.150 ;
        LAYER VTPH ;
        RECT  14.720 1.080 17.180 2.400 ;
        RECT  0.000 1.140 4.150 2.400 ;
        RECT  0.000 1.180 5.800 2.400 ;
        RECT  9.150 1.200 19.600 2.400 ;
        RECT  11.050 1.140 19.600 2.400 ;
        RECT  0.000 1.260 19.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 19.600 1.080 ;
        RECT  0.000 0.000 14.720 1.140 ;
        RECT  17.180 0.000 19.600 1.140 ;
        RECT  4.150 0.000 11.050 1.180 ;
        RECT  5.800 0.000 11.050 1.200 ;
        RECT  5.800 0.000 9.150 1.260 ;
    END
END SDFRM8HM

MACRO SDFRM4HM
    CLASS CORE ;
    FOREIGN SDFRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.481  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.010 2.860 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.190 1.050 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.583  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.900 1.380 15.410 1.600 ;
        RECT  14.900 0.470 15.410 0.670 ;
        RECT  14.900 0.470 15.120 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.330 1.440 17.100 1.640 ;
        RECT  16.900 0.660 17.100 1.640 ;
        RECT  16.330 0.660 17.100 0.860 ;
        RECT  16.330 1.440 16.530 2.080 ;
        RECT  16.330 0.430 16.530 0.860 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.293  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.700 1.120 13.440 1.280 ;
        RECT  11.700 0.840 12.000 1.280 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.200 2.540 ;
        RECT  16.850 1.840 17.050 2.540 ;
        RECT  15.730 2.080 16.010 2.540 ;
        RECT  14.520 2.080 14.800 2.540 ;
        RECT  13.500 1.770 13.780 2.540 ;
        RECT  12.460 1.760 12.740 2.540 ;
        RECT  11.540 1.500 11.700 2.540 ;
        RECT  11.420 1.500 11.700 1.700 ;
        RECT  8.700 2.080 8.980 2.540 ;
        RECT  4.360 2.020 4.560 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.200 0.140 ;
        RECT  16.810 -0.140 17.090 0.500 ;
        RECT  15.770 -0.140 15.970 0.650 ;
        RECT  14.580 -0.140 14.740 0.700 ;
        RECT  13.460 -0.140 13.740 0.320 ;
        RECT  11.020 -0.140 11.220 0.600 ;
        RECT  8.070 -0.140 8.350 0.710 ;
        RECT  4.660 -0.140 4.860 0.610 ;
        RECT  3.140 -0.140 3.420 0.500 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.700 ;
        RECT  0.140 1.540 1.640 1.700 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.900 0.620 4.180 1.300 ;
        RECT  3.720 1.100 4.770 1.300 ;
        RECT  3.720 1.100 3.880 1.760 ;
        RECT  4.040 1.700 4.880 1.860 ;
        RECT  2.600 1.760 3.520 1.920 ;
        RECT  1.620 1.860 1.910 2.100 ;
        RECT  3.360 1.760 3.520 2.100 ;
        RECT  4.720 1.700 4.880 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.040 1.700 4.200 2.100 ;
        RECT  3.360 1.940 4.200 2.100 ;
        RECT  5.520 1.740 5.720 2.100 ;
        RECT  4.720 1.940 5.720 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.580 0.300 4.500 0.460 ;
        RECT  5.020 0.300 6.060 0.460 ;
        RECT  5.860 0.300 6.060 0.600 ;
        RECT  2.820 0.300 2.980 0.820 ;
        RECT  1.840 0.300 2.000 0.690 ;
        RECT  4.340 0.300 4.500 0.930 ;
        RECT  3.580 0.300 3.740 0.820 ;
        RECT  2.820 0.660 3.740 0.820 ;
        RECT  5.020 0.300 5.180 0.930 ;
        RECT  4.340 0.770 5.180 0.930 ;
        RECT  6.220 0.300 7.100 0.460 ;
        RECT  6.900 0.300 7.100 0.700 ;
        RECT  5.340 0.660 5.620 0.920 ;
        RECT  6.220 0.300 6.380 0.920 ;
        RECT  5.340 0.760 6.380 0.920 ;
        RECT  5.340 0.660 5.540 1.450 ;
        RECT  5.040 1.250 5.540 1.450 ;
        RECT  5.040 1.250 5.240 1.780 ;
        RECT  6.780 1.620 8.220 1.780 ;
        RECT  6.540 0.980 8.320 1.140 ;
        RECT  6.540 0.620 6.740 1.240 ;
        RECT  6.040 1.080 6.740 1.240 ;
        RECT  6.040 1.080 6.240 2.020 ;
        RECT  8.800 0.600 9.000 1.600 ;
        RECT  7.160 1.300 9.000 1.460 ;
        RECT  8.800 1.440 9.660 1.600 ;
        RECT  9.460 1.440 9.660 1.780 ;
        RECT  8.380 1.760 9.300 1.920 ;
        RECT  9.140 1.760 9.300 2.100 ;
        RECT  8.380 1.760 8.540 2.100 ;
        RECT  6.400 1.940 8.540 2.100 ;
        RECT  9.140 1.940 9.820 2.100 ;
        RECT  9.440 0.300 10.340 0.460 ;
        RECT  10.180 0.300 10.340 1.420 ;
        RECT  9.440 0.300 9.640 1.280 ;
        RECT  10.180 1.220 10.760 1.420 ;
        RECT  9.820 0.620 10.020 1.780 ;
        RECT  9.820 1.620 10.660 1.780 ;
        RECT  10.490 1.620 10.660 2.100 ;
        RECT  10.490 1.940 11.360 2.100 ;
        RECT  12.460 0.620 12.740 0.960 ;
        RECT  12.460 0.800 14.080 0.960 ;
        RECT  13.880 0.800 14.080 1.600 ;
        RECT  12.000 1.440 14.080 1.600 ;
        RECT  12.000 1.440 12.160 1.840 ;
        RECT  13.020 1.440 13.220 1.870 ;
        RECT  11.380 0.300 13.190 0.460 ;
        RECT  13.030 0.300 13.190 0.640 ;
        RECT  13.030 0.480 14.400 0.640 ;
        RECT  10.500 0.480 10.700 1.000 ;
        RECT  11.380 0.300 11.540 1.000 ;
        RECT  10.500 0.840 11.540 1.000 ;
        RECT  15.650 1.040 16.550 1.240 ;
        RECT  14.240 0.480 14.400 1.920 ;
        RECT  10.980 0.840 11.180 1.780 ;
        RECT  15.650 1.040 15.850 1.920 ;
        RECT  13.980 1.760 15.850 1.920 ;
        LAYER VI1 ;
        RECT  6.900 0.380 7.100 0.580 ;
        RECT  9.440 0.850 9.640 1.050 ;
        LAYER ME2 ;
        RECT  6.750 0.380 9.640 0.580 ;
        RECT  9.440 0.380 9.640 1.150 ;
        LAYER VTPH ;
        RECT  14.570 1.080 15.750 2.400 ;
        RECT  0.000 1.140 4.150 2.400 ;
        RECT  0.000 1.200 5.800 2.400 ;
        RECT  9.220 1.200 17.200 2.400 ;
        RECT  10.350 1.140 17.200 2.400 ;
        RECT  0.000 1.260 17.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.200 1.080 ;
        RECT  0.000 0.000 14.570 1.140 ;
        RECT  15.750 0.000 17.200 1.140 ;
        RECT  4.150 0.000 10.350 1.200 ;
        RECT  5.800 0.000 9.220 1.260 ;
    END
END SDFRM4HM

MACRO SDFRM2HM
    CLASS CORE ;
    FOREIGN SDFRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.481  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.010 2.860 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.190 1.050 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.980 1.380 14.300 1.600 ;
        RECT  14.060 0.470 14.300 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.180 1.440 15.500 2.080 ;
        RECT  15.300 0.470 15.500 2.080 ;
        RECT  15.140 0.470 15.500 0.670 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.700 0.840 12.040 1.250 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  14.580 2.080 14.860 2.540 ;
        RECT  13.420 2.080 13.700 2.540 ;
        RECT  12.460 1.730 12.740 2.540 ;
        RECT  11.540 1.500 11.700 2.540 ;
        RECT  11.420 1.500 11.700 1.700 ;
        RECT  8.700 2.080 8.980 2.540 ;
        RECT  4.360 2.020 4.560 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  14.580 -0.140 14.780 0.760 ;
        RECT  13.580 -0.140 13.780 0.750 ;
        RECT  11.020 -0.140 11.220 0.600 ;
        RECT  8.070 -0.140 8.350 0.710 ;
        RECT  4.660 -0.140 4.860 0.610 ;
        RECT  3.140 -0.140 3.420 0.500 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.700 ;
        RECT  0.140 1.540 1.640 1.700 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.900 0.620 4.180 1.300 ;
        RECT  3.720 1.100 4.770 1.300 ;
        RECT  3.720 1.100 3.880 1.760 ;
        RECT  4.040 1.700 4.880 1.860 ;
        RECT  2.600 1.760 3.520 1.920 ;
        RECT  1.620 1.860 1.910 2.100 ;
        RECT  3.360 1.760 3.520 2.100 ;
        RECT  4.720 1.700 4.880 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.040 1.700 4.200 2.100 ;
        RECT  3.360 1.940 4.200 2.100 ;
        RECT  5.520 1.740 5.720 2.100 ;
        RECT  4.720 1.940 5.720 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.580 0.300 4.500 0.460 ;
        RECT  5.020 0.300 6.060 0.460 ;
        RECT  5.860 0.300 6.060 0.600 ;
        RECT  2.820 0.300 2.980 0.820 ;
        RECT  1.840 0.300 2.000 0.690 ;
        RECT  4.340 0.300 4.500 0.930 ;
        RECT  3.580 0.300 3.740 0.820 ;
        RECT  2.820 0.660 3.740 0.820 ;
        RECT  5.020 0.300 5.180 0.930 ;
        RECT  4.340 0.770 5.180 0.930 ;
        RECT  6.220 0.300 7.100 0.460 ;
        RECT  6.900 0.300 7.100 0.700 ;
        RECT  5.340 0.660 5.620 0.920 ;
        RECT  6.220 0.300 6.380 0.920 ;
        RECT  5.340 0.760 6.380 0.920 ;
        RECT  5.340 0.660 5.540 1.450 ;
        RECT  5.040 1.250 5.540 1.450 ;
        RECT  5.040 1.250 5.240 1.780 ;
        RECT  6.640 1.500 6.840 1.780 ;
        RECT  6.640 1.620 8.220 1.780 ;
        RECT  6.540 0.980 8.320 1.140 ;
        RECT  6.540 0.620 6.740 1.240 ;
        RECT  6.040 1.080 6.740 1.240 ;
        RECT  6.040 1.080 6.240 2.020 ;
        RECT  8.800 0.600 9.000 1.600 ;
        RECT  7.000 1.300 9.000 1.460 ;
        RECT  8.800 1.440 9.660 1.600 ;
        RECT  9.460 1.440 9.660 1.780 ;
        RECT  8.380 1.760 9.300 1.920 ;
        RECT  9.140 1.760 9.300 2.100 ;
        RECT  8.380 1.760 8.540 2.100 ;
        RECT  6.400 1.940 8.540 2.100 ;
        RECT  9.140 1.940 9.820 2.100 ;
        RECT  9.440 0.300 10.340 0.460 ;
        RECT  10.180 0.300 10.340 1.420 ;
        RECT  9.440 0.300 9.640 1.280 ;
        RECT  10.180 1.220 10.760 1.420 ;
        RECT  9.820 0.620 10.020 1.780 ;
        RECT  9.820 1.620 10.660 1.780 ;
        RECT  10.490 1.620 10.660 2.100 ;
        RECT  10.490 1.940 11.360 2.100 ;
        RECT  12.460 0.620 12.740 1.240 ;
        RECT  12.460 0.960 12.840 1.240 ;
        RECT  12.460 0.620 12.690 1.570 ;
        RECT  11.980 1.410 12.690 1.570 ;
        RECT  11.980 1.410 12.180 1.770 ;
        RECT  11.380 0.300 13.160 0.460 ;
        RECT  10.500 0.480 10.700 1.000 ;
        RECT  11.380 0.300 11.540 1.000 ;
        RECT  10.500 0.840 11.540 1.000 ;
        RECT  14.460 1.040 15.080 1.240 ;
        RECT  13.000 0.300 13.160 1.920 ;
        RECT  10.980 0.840 11.180 1.780 ;
        RECT  14.460 1.040 14.660 1.920 ;
        RECT  13.000 1.760 14.660 1.920 ;
        LAYER VI1 ;
        RECT  6.900 0.380 7.100 0.580 ;
        RECT  9.440 0.850 9.640 1.050 ;
        LAYER ME2 ;
        RECT  6.750 0.380 9.640 0.580 ;
        RECT  9.440 0.380 9.640 1.150 ;
        LAYER VTPH ;
        RECT  12.960 1.080 14.800 2.400 ;
        RECT  0.000 1.140 4.150 2.400 ;
        RECT  0.000 1.200 7.440 2.400 ;
        RECT  9.220 1.200 15.600 2.400 ;
        RECT  10.350 1.140 15.600 2.400 ;
        RECT  0.000 1.260 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.080 ;
        RECT  0.000 0.000 12.960 1.140 ;
        RECT  14.800 0.000 15.600 1.140 ;
        RECT  4.150 0.000 10.350 1.200 ;
        RECT  7.440 0.000 9.220 1.260 ;
    END
END SDFRM2HM

MACRO SDFRM1HM
    CLASS CORE ;
    FOREIGN SDFRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.438  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.920 0.990 2.120 1.190 ;
        LAYER ME2 ;
        RECT  1.830 0.840 2.300 1.220 ;
        LAYER ME1 ;
        RECT  1.880 0.930 2.160 1.380 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.840 3.290 1.280 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.340  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.700 0.470 14.020 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.900 0.430 15.140 1.860 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.520 0.840 11.900 1.250 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.870 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  14.340 2.080 14.620 2.540 ;
        RECT  13.180 2.080 13.460 2.540 ;
        RECT  12.220 1.730 12.500 2.540 ;
        RECT  11.300 1.500 11.460 2.540 ;
        RECT  11.180 1.500 11.460 1.700 ;
        RECT  8.460 2.080 8.740 2.540 ;
        RECT  4.300 2.020 4.500 2.540 ;
        RECT  2.960 1.800 3.180 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  14.340 -0.140 14.540 0.760 ;
        RECT  13.340 -0.140 13.540 0.750 ;
        RECT  10.780 -0.140 10.980 0.600 ;
        RECT  7.660 -0.140 7.940 0.540 ;
        RECT  4.300 -0.140 4.500 0.610 ;
        RECT  2.660 -0.140 2.940 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.500 0.810 2.660 1.280 ;
        RECT  2.320 1.120 2.660 1.280 ;
        RECT  1.440 1.070 1.640 1.700 ;
        RECT  2.320 1.120 2.480 1.700 ;
        RECT  0.140 1.540 2.480 1.700 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  3.540 0.620 3.820 0.840 ;
        RECT  3.660 1.100 4.710 1.300 ;
        RECT  3.660 0.620 3.820 1.760 ;
        RECT  2.640 1.480 3.500 1.640 ;
        RECT  3.980 1.700 4.820 1.860 ;
        RECT  3.340 1.480 3.500 2.100 ;
        RECT  4.660 1.700 4.820 2.100 ;
        RECT  2.640 1.480 2.800 2.020 ;
        RECT  1.580 1.860 2.800 2.020 ;
        RECT  3.980 1.700 4.140 2.100 ;
        RECT  3.340 1.940 4.140 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.660 1.940 5.660 2.100 ;
        RECT  3.100 0.300 4.140 0.460 ;
        RECT  4.660 0.300 5.700 0.460 ;
        RECT  1.820 0.370 2.020 0.650 ;
        RECT  5.500 0.300 5.700 0.600 ;
        RECT  3.100 0.300 3.260 0.650 ;
        RECT  1.820 0.490 3.260 0.650 ;
        RECT  3.980 0.300 4.140 0.930 ;
        RECT  4.660 0.300 4.820 0.930 ;
        RECT  3.980 0.770 4.820 0.930 ;
        RECT  5.860 0.300 6.820 0.460 ;
        RECT  6.620 0.300 6.820 0.700 ;
        RECT  4.980 0.660 5.260 0.920 ;
        RECT  5.860 0.300 6.020 0.920 ;
        RECT  4.980 0.760 6.020 0.920 ;
        RECT  4.980 0.660 5.180 1.780 ;
        RECT  6.580 1.500 6.780 1.780 ;
        RECT  6.580 1.620 7.980 1.780 ;
        RECT  6.180 0.680 6.460 1.340 ;
        RECT  5.980 1.180 8.000 1.340 ;
        RECT  7.800 1.180 8.000 1.460 ;
        RECT  5.980 1.180 6.180 2.020 ;
        RECT  7.000 0.300 7.200 0.860 ;
        RECT  7.000 0.700 8.460 0.860 ;
        RECT  8.260 0.600 8.460 1.600 ;
        RECT  8.260 1.440 9.420 1.600 ;
        RECT  9.220 1.440 9.420 1.780 ;
        RECT  8.140 1.760 9.060 1.920 ;
        RECT  8.900 1.760 9.060 2.100 ;
        RECT  8.140 1.760 8.300 2.100 ;
        RECT  6.340 1.940 8.300 2.100 ;
        RECT  8.900 1.940 9.580 2.100 ;
        RECT  8.980 0.300 10.100 0.460 ;
        RECT  9.940 0.300 10.100 1.420 ;
        RECT  8.980 0.300 9.180 1.230 ;
        RECT  9.940 1.220 10.520 1.420 ;
        RECT  9.580 0.620 9.780 1.780 ;
        RECT  9.580 1.620 10.420 1.780 ;
        RECT  10.250 1.620 10.420 2.100 ;
        RECT  10.250 1.940 11.120 2.100 ;
        RECT  12.220 0.620 12.500 1.240 ;
        RECT  12.220 0.960 12.600 1.240 ;
        RECT  12.220 0.620 12.450 1.570 ;
        RECT  11.740 1.410 12.450 1.570 ;
        RECT  11.740 1.410 11.940 1.770 ;
        RECT  11.140 0.300 12.920 0.460 ;
        RECT  10.260 0.480 10.460 1.000 ;
        RECT  11.140 0.300 11.300 1.000 ;
        RECT  10.260 0.840 11.300 1.000 ;
        RECT  14.220 1.040 14.720 1.240 ;
        RECT  12.760 0.300 12.920 1.920 ;
        RECT  10.740 0.840 10.940 1.780 ;
        RECT  14.220 1.040 14.420 1.920 ;
        RECT  12.760 1.760 14.420 1.920 ;
        LAYER VI1 ;
        RECT  6.620 0.380 6.820 0.580 ;
        RECT  8.980 0.800 9.180 1.000 ;
        LAYER ME2 ;
        RECT  6.520 0.380 9.180 0.580 ;
        RECT  8.980 0.380 9.180 1.100 ;
        LAYER VTPH ;
        RECT  1.520 1.050 2.600 2.400 ;
        RECT  12.720 1.080 14.560 2.400 ;
        RECT  0.000 1.140 4.100 2.400 ;
        RECT  0.000 1.200 7.000 2.400 ;
        RECT  8.680 1.200 15.600 2.400 ;
        RECT  10.110 1.140 15.600 2.400 ;
        RECT  0.000 1.260 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.050 ;
        RECT  2.600 0.000 15.600 1.080 ;
        RECT  0.000 0.000 1.520 1.140 ;
        RECT  2.600 0.000 12.720 1.140 ;
        RECT  14.560 0.000 15.600 1.140 ;
        RECT  4.100 0.000 10.110 1.200 ;
        RECT  7.000 0.000 8.680 1.260 ;
    END
END SDFRM1HM

MACRO SDFQZRM8HM
    CLASS CORE ;
    FOREIGN SDFQZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.312  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.320 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        ANTENNAGATEAREA 0.146  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.628  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.070 0.430 16.400 2.100 ;
        RECT  14.890 0.900 16.400 1.100 ;
        RECT  15.100 0.430 15.300 1.100 ;
        RECT  14.890 0.900 15.190 2.100 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.570 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.200 2.540 ;
        RECT  16.660 1.480 16.860 2.540 ;
        RECT  15.620 1.420 15.820 2.540 ;
        RECT  14.260 1.840 14.460 2.540 ;
        RECT  12.980 1.840 13.260 2.540 ;
        RECT  10.600 1.800 10.760 2.540 ;
        RECT  9.160 2.080 9.440 2.540 ;
        RECT  5.820 1.840 6.020 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.200 0.140 ;
        RECT  16.670 -0.140 16.870 0.710 ;
        RECT  15.620 -0.140 15.820 0.710 ;
        RECT  14.580 -0.140 14.780 0.710 ;
        RECT  13.600 -0.140 13.760 0.700 ;
        RECT  10.600 -0.140 10.880 0.500 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.380 1.420 0.580 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.380 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.340 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  6.780 0.620 7.060 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.500 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.300 0.300 7.500 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  8.040 0.620 8.240 1.080 ;
        RECT  8.040 0.880 9.620 1.080 ;
        RECT  8.040 0.620 8.220 1.740 ;
        RECT  8.040 1.540 8.420 1.740 ;
        RECT  8.880 1.240 9.080 1.600 ;
        RECT  9.840 0.620 10.120 1.600 ;
        RECT  8.880 1.440 10.120 1.600 ;
        RECT  9.920 0.620 10.120 1.780 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.340 0.960 ;
        RECT  10.280 1.360 10.920 1.560 ;
        RECT  5.300 1.480 6.340 1.680 ;
        RECT  5.300 1.480 5.500 1.920 ;
        RECT  8.840 1.760 9.760 1.920 ;
        RECT  6.180 0.800 6.340 2.100 ;
        RECT  9.600 1.760 9.760 2.100 ;
        RECT  8.840 1.760 9.000 2.100 ;
        RECT  6.180 1.940 9.000 2.100 ;
        RECT  10.280 1.360 10.440 2.100 ;
        RECT  9.600 1.940 10.440 2.100 ;
        RECT  11.040 0.300 11.540 0.600 ;
        RECT  7.680 0.300 8.560 0.460 ;
        RECT  9.360 0.300 10.440 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  9.360 0.300 9.520 0.720 ;
        RECT  8.400 0.560 9.520 0.720 ;
        RECT  10.280 0.300 10.440 0.980 ;
        RECT  10.280 0.780 11.600 0.980 ;
        RECT  11.380 0.780 11.600 1.100 ;
        RECT  7.680 0.300 7.880 1.540 ;
        RECT  11.760 0.300 11.960 1.700 ;
        RECT  11.490 1.540 11.960 1.700 ;
        RECT  12.660 0.620 13.120 0.900 ;
        RECT  12.300 0.300 13.440 0.460 ;
        RECT  12.300 0.300 12.500 0.700 ;
        RECT  13.280 0.300 13.440 1.280 ;
        RECT  12.120 1.080 13.840 1.280 ;
        RECT  12.120 1.080 12.280 2.020 ;
        RECT  10.980 1.860 12.280 2.020 ;
        RECT  14.100 0.430 14.300 1.680 ;
        RECT  12.760 1.480 14.300 1.680 ;
        LAYER VI1 ;
        RECT  6.780 1.200 6.980 1.400 ;
        RECT  7.680 1.200 7.880 1.400 ;
        RECT  9.920 0.960 10.120 1.160 ;
        RECT  10.620 1.360 10.820 1.560 ;
        RECT  11.140 0.400 11.340 0.600 ;
        RECT  11.760 0.960 11.960 1.160 ;
        RECT  12.300 0.400 12.500 0.600 ;
        RECT  12.820 0.620 13.020 0.820 ;
        LAYER ME2 ;
        RECT  6.680 1.200 7.980 1.400 ;
        RECT  9.840 0.960 12.020 1.160 ;
        RECT  11.040 0.400 12.600 0.600 ;
        RECT  12.820 0.520 13.020 1.560 ;
        RECT  10.520 1.360 13.020 1.560 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  10.810 1.090 12.520 2.400 ;
        RECT  0.000 1.140 7.770 2.400 ;
        RECT  8.800 1.140 17.200 2.400 ;
        RECT  0.000 1.200 17.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.200 1.080 ;
        RECT  4.080 0.000 17.200 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 10.810 1.140 ;
        RECT  12.520 0.000 17.200 1.140 ;
        RECT  7.770 0.000 8.800 1.200 ;
    END
END SDFQZRM8HM

MACRO SDFQZRM4HM
    CLASS CORE ;
    FOREIGN SDFQZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        ANTENNAGATEAREA 0.078  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.933  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.312  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.380 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.340 0.390 13.660 2.100 ;
        RECT  13.200 0.840 13.660 1.160 ;
        RECT  13.330 0.390 13.660 1.160 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.570 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.400 2.540 ;
        RECT  13.920 1.400 14.120 2.540 ;
        RECT  12.840 1.400 13.040 2.540 ;
        RECT  11.630 1.840 11.910 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.820 1.840 6.020 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.400 0.140 ;
        RECT  13.930 -0.140 14.130 0.670 ;
        RECT  12.890 -0.140 13.090 0.670 ;
        RECT  11.910 -0.140 12.070 0.700 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.380 1.420 0.580 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.380 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.340 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  6.780 0.620 7.060 1.400 ;
        RECT  6.540 1.220 7.060 1.400 ;
        RECT  6.540 1.220 6.740 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.480 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.220 0.300 7.480 0.660 ;
        RECT  7.220 0.300 7.380 1.780 ;
        RECT  6.980 1.580 7.380 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  7.960 0.880 9.460 1.080 ;
        RECT  7.960 0.620 8.160 1.780 ;
        RECT  7.880 1.580 8.160 1.780 ;
        RECT  7.640 0.300 8.560 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  8.400 0.560 9.880 0.720 ;
        RECT  7.640 0.300 7.800 1.000 ;
        RECT  9.720 0.560 9.880 1.090 ;
        RECT  7.540 0.850 7.700 1.490 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.340 0.960 ;
        RECT  5.300 1.500 6.340 1.680 ;
        RECT  8.420 1.720 9.560 1.920 ;
        RECT  6.180 0.800 6.340 2.100 ;
        RECT  5.300 1.500 5.500 2.050 ;
        RECT  8.420 1.720 8.580 2.100 ;
        RECT  6.180 1.940 8.580 2.100 ;
        RECT  9.400 1.900 10.080 2.100 ;
        RECT  10.040 0.300 10.200 1.460 ;
        RECT  8.700 1.300 10.200 1.460 ;
        RECT  9.720 1.300 9.920 1.720 ;
        RECT  10.940 0.620 11.400 0.900 ;
        RECT  10.560 0.300 11.720 0.460 ;
        RECT  10.560 0.300 10.760 0.660 ;
        RECT  11.560 0.300 11.720 1.280 ;
        RECT  10.580 1.080 12.120 1.280 ;
        RECT  10.580 1.080 10.740 1.950 ;
        RECT  12.410 0.390 12.610 1.680 ;
        RECT  11.220 1.480 12.610 1.680 ;
        LAYER VI1 ;
        RECT  9.200 1.720 9.400 1.920 ;
        RECT  11.100 0.620 11.300 0.820 ;
        LAYER ME2 ;
        RECT  11.100 0.520 11.300 1.920 ;
        RECT  9.100 1.720 11.300 1.920 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  8.800 1.090 10.980 2.400 ;
        RECT  0.000 1.140 5.840 2.400 ;
        RECT  8.800 1.140 14.400 2.400 ;
        RECT  0.000 1.200 14.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.400 1.080 ;
        RECT  4.080 0.000 14.400 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 8.800 1.140 ;
        RECT  10.980 0.000 14.400 1.140 ;
        RECT  5.840 0.000 8.800 1.200 ;
    END
END SDFQZRM4HM

MACRO SDFQZRM2HM
    CLASS CORE ;
    FOREIGN SDFQZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        ANTENNAGATEAREA 0.078  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.933  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.312  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.320 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.900 0.390 13.100 1.160 ;
        RECT  12.740 0.950 13.000 2.100 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.570 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.260 1.400 13.460 2.540 ;
        RECT  11.640 1.840 11.840 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.820 1.840 6.020 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.420 -0.140 13.620 0.670 ;
        RECT  11.780 -0.140 11.940 0.610 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.380 1.420 0.580 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.380 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.340 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  6.780 0.620 7.060 1.400 ;
        RECT  6.540 1.220 7.060 1.400 ;
        RECT  6.540 1.220 6.740 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.480 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.220 0.300 7.480 0.660 ;
        RECT  7.220 0.300 7.380 1.780 ;
        RECT  6.980 1.580 7.380 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  7.960 0.880 9.460 1.080 ;
        RECT  7.960 0.620 8.160 1.780 ;
        RECT  7.880 1.580 8.160 1.780 ;
        RECT  7.640 0.300 8.560 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  8.400 0.560 9.880 0.720 ;
        RECT  7.640 0.300 7.800 1.000 ;
        RECT  9.720 0.560 9.880 1.090 ;
        RECT  7.540 0.850 7.700 1.490 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.340 0.960 ;
        RECT  5.300 1.500 6.340 1.680 ;
        RECT  8.420 1.720 9.560 1.920 ;
        RECT  6.180 0.800 6.340 2.100 ;
        RECT  5.300 1.500 5.500 2.050 ;
        RECT  8.420 1.720 8.580 2.100 ;
        RECT  6.180 1.940 8.580 2.100 ;
        RECT  9.400 1.900 10.080 2.100 ;
        RECT  10.040 0.300 10.200 1.460 ;
        RECT  8.700 1.300 10.200 1.460 ;
        RECT  9.720 1.300 9.920 1.720 ;
        RECT  10.920 0.620 11.380 0.900 ;
        RECT  12.060 1.000 12.260 1.280 ;
        RECT  10.560 1.080 12.260 1.280 ;
        RECT  10.560 0.380 10.760 2.070 ;
        RECT  12.320 0.300 12.580 0.580 ;
        RECT  12.420 0.300 12.580 1.680 ;
        RECT  11.220 1.480 12.580 1.680 ;
        LAYER VI1 ;
        RECT  9.200 1.720 9.400 1.920 ;
        RECT  11.080 0.620 11.280 0.820 ;
        LAYER ME2 ;
        RECT  11.080 0.520 11.280 1.920 ;
        RECT  9.100 1.720 11.280 1.920 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  8.800 1.090 10.980 2.400 ;
        RECT  0.000 1.140 5.840 2.400 ;
        RECT  8.800 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  4.080 0.000 14.000 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 8.800 1.140 ;
        RECT  10.980 0.000 14.000 1.140 ;
        RECT  5.840 0.000 8.800 1.200 ;
    END
END SDFQZRM2HM

MACRO SDFQZRM1HM
    CLASS CORE ;
    FOREIGN SDFQZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        ANTENNAGATEAREA 0.053  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.288  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.120 5.500 1.320 ;
        LAYER ME2 ;
        RECT  5.300 1.020 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.180 1.120 5.720 1.320 ;
        END
    END CK
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        ANTENNAGATEAREA 0.065  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.099  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.020 3.100 1.220 ;
        LAYER ME2 ;
        RECT  2.850 0.750 3.100 1.320 ;
        LAYER ME1 ;
        RECT  2.720 1.020 3.220 1.280 ;
        END
    END SD
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.730 0.840 13.150 1.160 ;
        RECT  12.730 0.390 13.020 1.160 ;
        RECT  12.730 0.390 12.990 2.010 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.250 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 0.700 3.540 1.280 ;
        RECT  1.900 0.700 3.540 0.860 ;
        RECT  1.900 0.440 2.300 0.860 ;
        RECT  1.900 0.440 2.060 1.600 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.290 1.770 13.490 2.540 ;
        RECT  11.690 1.840 11.890 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.900 1.840 6.100 2.540 ;
        RECT  4.220 2.080 4.500 2.540 ;
        RECT  3.020 2.080 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.290 -0.140 13.490 0.670 ;
        RECT  11.710 -0.140 11.870 0.610 ;
        RECT  9.000 -0.140 9.200 0.390 ;
        RECT  6.020 -0.140 6.300 0.320 ;
        RECT  4.300 -0.140 4.500 0.710 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  0.140 -0.140 0.340 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.940 0.400 1.420 0.600 ;
        RECT  0.140 1.460 1.420 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.260 0.400 1.420 2.100 ;
        RECT  1.180 1.460 1.420 2.100 ;
        RECT  3.580 0.380 3.940 0.540 ;
        RECT  2.360 1.260 2.560 1.600 ;
        RECT  3.780 0.380 3.940 1.600 ;
        RECT  2.360 1.440 3.940 1.600 ;
        RECT  1.580 0.320 1.740 1.920 ;
        RECT  4.360 1.020 4.560 1.920 ;
        RECT  1.580 1.760 4.560 1.920 ;
        RECT  1.880 1.760 2.080 2.100 ;
        RECT  6.780 0.620 7.060 1.400 ;
        RECT  6.580 1.220 6.780 1.780 ;
        RECT  4.820 0.300 5.860 0.460 ;
        RECT  6.460 0.300 7.480 0.460 ;
        RECT  5.700 0.300 5.860 0.640 ;
        RECT  6.460 0.300 6.620 0.640 ;
        RECT  5.700 0.480 6.620 0.640 ;
        RECT  7.220 0.300 7.480 0.660 ;
        RECT  7.220 0.300 7.380 1.780 ;
        RECT  7.020 1.580 7.380 1.780 ;
        RECT  4.820 0.300 5.020 2.100 ;
        RECT  7.960 0.880 9.460 1.080 ;
        RECT  7.960 0.620 8.160 1.780 ;
        RECT  7.880 1.580 8.160 1.780 ;
        RECT  7.640 0.300 8.560 0.460 ;
        RECT  8.400 0.300 8.560 0.720 ;
        RECT  8.400 0.560 9.880 0.720 ;
        RECT  7.640 0.300 7.800 1.000 ;
        RECT  9.720 0.560 9.880 1.090 ;
        RECT  7.540 0.850 7.700 1.490 ;
        RECT  5.260 0.620 5.540 0.960 ;
        RECT  5.260 0.800 6.420 0.960 ;
        RECT  5.300 1.500 6.420 1.680 ;
        RECT  8.420 1.720 9.560 1.920 ;
        RECT  6.260 0.800 6.420 2.100 ;
        RECT  5.300 1.500 5.500 2.100 ;
        RECT  8.420 1.720 8.580 2.100 ;
        RECT  6.260 1.940 8.580 2.100 ;
        RECT  9.400 1.900 10.080 2.100 ;
        RECT  10.040 0.300 10.200 1.460 ;
        RECT  8.700 1.300 10.200 1.460 ;
        RECT  9.720 1.300 9.920 1.720 ;
        RECT  10.970 0.510 11.430 0.900 ;
        RECT  11.750 1.000 12.100 1.280 ;
        RECT  10.560 1.080 12.100 1.280 ;
        RECT  10.560 0.380 10.760 2.070 ;
        RECT  12.250 0.300 12.510 0.580 ;
        RECT  12.260 0.300 12.510 1.680 ;
        RECT  11.270 1.480 12.510 1.680 ;
        RECT  12.280 0.300 12.510 1.800 ;
        LAYER VI1 ;
        RECT  9.100 1.720 9.300 1.920 ;
        RECT  11.010 0.620 11.210 0.820 ;
        LAYER ME2 ;
        RECT  10.970 0.520 11.210 1.920 ;
        RECT  9.000 1.720 11.210 1.920 ;
        LAYER VTPH ;
        RECT  3.440 1.080 4.080 2.400 ;
        RECT  8.800 1.090 11.030 2.400 ;
        RECT  0.000 1.140 5.840 2.400 ;
        RECT  8.800 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  4.080 0.000 14.000 1.090 ;
        RECT  0.000 0.000 3.440 1.140 ;
        RECT  4.080 0.000 8.800 1.140 ;
        RECT  11.030 0.000 14.000 1.140 ;
        RECT  5.840 0.000 8.800 1.200 ;
    END
END SDFQZRM1HM

MACRO SDFQSM8HM
    CLASS CORE ;
    FOREIGN SDFQSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.220 0.840 7.500 1.250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.620 3.240 3.100 3.700 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.440 1.900 2.080 ;
        RECT  0.900 0.660 1.900 0.860 ;
        RECT  1.700 0.440 1.900 0.860 ;
        RECT  0.660 1.440 1.900 1.640 ;
        RECT  0.900 0.660 1.100 1.640 ;
        RECT  0.660 0.660 1.900 0.830 ;
        RECT  0.660 1.440 0.860 2.080 ;
        RECT  0.660 0.440 0.860 0.830 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.000 1.120 4.300 1.560 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 3.550 1.160 4.000 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.550 0.700 4.100 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.420 1.540 7.620 3.260 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.780 2.260 3.060 2.640 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.660 2.260 0.940 2.960 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.420 -0.140 7.620 0.660 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.710 ;
        RECT  0.000 4.660 8.000 4.940 ;
        RECT  7.420 4.180 7.620 4.940 ;
        RECT  4.700 4.480 4.980 4.940 ;
        RECT  2.940 4.240 3.140 4.940 ;
        RECT  0.660 4.260 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.120 1.500 3.280 ;
        RECT  1.340 3.120 1.500 3.850 ;
        RECT  1.340 3.650 2.000 3.850 ;
        RECT  0.140 3.030 0.340 4.270 ;
        RECT  2.180 3.120 2.460 4.180 ;
        RECT  2.740 0.440 2.940 0.860 ;
        RECT  2.220 0.660 2.940 0.860 ;
        RECT  1.480 1.040 2.420 1.240 ;
        RECT  2.220 0.660 2.420 1.570 ;
        RECT  3.480 1.060 3.680 1.570 ;
        RECT  2.220 1.380 3.680 1.570 ;
        RECT  2.740 1.380 2.940 2.080 ;
        RECT  3.940 3.780 4.600 4.000 ;
        RECT  3.940 3.780 4.220 4.180 ;
        RECT  4.090 0.640 4.620 0.800 ;
        RECT  4.460 1.750 5.180 1.950 ;
        RECT  4.460 0.640 4.620 2.050 ;
        RECT  3.820 1.850 4.620 2.050 ;
        RECT  3.700 0.320 5.120 0.480 ;
        RECT  3.700 0.320 3.860 0.820 ;
        RECT  3.100 0.660 3.860 0.820 ;
        RECT  3.100 0.660 3.260 1.220 ;
        RECT  2.700 1.060 3.260 1.220 ;
        RECT  4.960 0.320 5.120 1.520 ;
        RECT  4.960 1.360 5.900 1.520 ;
        RECT  5.700 1.360 5.900 1.900 ;
        RECT  3.280 3.440 5.080 3.600 ;
        RECT  3.280 3.440 3.480 3.760 ;
        RECT  4.800 3.360 5.080 4.000 ;
        RECT  4.800 3.840 5.940 4.000 ;
        RECT  5.660 3.840 5.940 4.180 ;
        RECT  3.280 2.720 6.140 2.880 ;
        RECT  1.660 2.800 3.420 2.960 ;
        RECT  1.660 2.800 1.860 3.080 ;
        RECT  2.620 3.920 3.460 4.080 ;
        RECT  4.380 4.160 5.300 4.320 ;
        RECT  1.660 4.140 1.860 4.500 ;
        RECT  3.300 3.920 3.460 4.500 ;
        RECT  5.140 4.160 5.300 4.500 ;
        RECT  2.620 3.920 2.780 4.500 ;
        RECT  1.660 4.340 2.780 4.500 ;
        RECT  4.380 4.160 4.540 4.500 ;
        RECT  3.300 4.340 4.540 4.500 ;
        RECT  6.220 4.050 6.420 4.500 ;
        RECT  5.140 4.340 6.420 4.500 ;
        RECT  5.460 0.600 5.660 1.200 ;
        RECT  5.460 1.040 6.450 1.200 ;
        RECT  6.250 1.040 6.450 1.900 ;
        RECT  6.300 2.700 6.740 2.860 ;
        RECT  4.320 3.040 6.460 3.200 ;
        RECT  6.300 2.700 6.460 3.200 ;
        RECT  3.380 3.120 4.600 3.280 ;
        RECT  5.360 3.480 7.060 3.640 ;
        RECT  6.860 3.080 7.060 4.330 ;
        RECT  5.840 0.380 7.060 0.580 ;
        RECT  6.860 0.380 7.060 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.550 3.660 ;
        RECT  6.490 1.140 8.000 3.660 ;
        RECT  0.000 1.180 8.000 3.660 ;
        RECT  4.510 1.180 5.370 3.880 ;
        LAYER VTNH ;
        RECT  0.000 3.660 4.510 4.800 ;
        RECT  5.370 3.660 8.000 4.800 ;
        RECT  0.000 3.880 8.000 4.800 ;
        RECT  0.000 0.000 8.000 1.140 ;
        RECT  3.550 0.000 6.490 1.180 ;
    END
END SDFQSM8HM

MACRO SDFQSM4HM
    CLASS CORE ;
    FOREIGN SDFQSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.411  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.530 1.080 2.730 1.280 ;
        LAYER ME2 ;
        RECT  2.500 0.950 2.760 1.450 ;
        LAYER ME1 ;
        RECT  2.460 1.050 2.900 1.300 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.200 1.020 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.880 1.440 14.300 1.640 ;
        RECT  14.100 0.710 14.300 1.640 ;
        RECT  13.880 0.710 14.300 0.870 ;
        RECT  13.880 1.440 14.080 2.080 ;
        RECT  13.880 0.450 14.080 0.870 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.900 1.200 11.200 1.590 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.750 1.140 1.250 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 0.720 1.250 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  14.400 1.840 14.600 2.540 ;
        RECT  13.360 1.840 13.560 2.540 ;
        RECT  12.300 1.840 12.500 2.540 ;
        RECT  11.060 2.080 11.340 2.540 ;
        RECT  8.550 1.830 8.840 2.540 ;
        RECT  7.030 2.080 7.310 2.540 ;
        RECT  4.300 1.980 4.460 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  14.400 -0.140 14.600 0.570 ;
        RECT  13.320 -0.140 13.600 0.500 ;
        RECT  12.280 -0.140 12.560 0.500 ;
        RECT  11.690 -0.140 11.970 0.500 ;
        RECT  7.230 -0.140 7.510 0.320 ;
        RECT  4.510 -0.140 4.670 0.420 ;
        RECT  3.060 -0.140 3.260 0.380 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 1.050 1.620 1.700 ;
        RECT  0.140 1.540 1.620 1.700 ;
        RECT  0.140 0.530 0.340 1.750 ;
        RECT  2.140 0.620 2.580 0.840 ;
        RECT  2.140 0.620 2.300 1.690 ;
        RECT  2.140 1.470 2.420 1.690 ;
        RECT  3.740 0.620 4.020 1.210 ;
        RECT  3.660 1.010 4.620 1.210 ;
        RECT  3.660 1.010 3.820 1.760 ;
        RECT  3.980 1.660 4.800 1.820 ;
        RECT  2.580 1.760 3.500 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  4.640 1.660 4.800 2.100 ;
        RECT  2.580 1.760 2.740 2.100 ;
        RECT  1.620 1.940 2.740 2.100 ;
        RECT  3.980 1.660 4.140 2.100 ;
        RECT  3.340 1.940 4.140 2.100 ;
        RECT  5.470 1.640 5.670 2.100 ;
        RECT  4.640 1.940 5.670 2.100 ;
        RECT  1.780 0.300 2.900 0.460 ;
        RECT  3.420 0.300 4.340 0.460 ;
        RECT  4.850 0.330 5.870 0.490 ;
        RECT  2.740 0.300 2.900 0.700 ;
        RECT  4.180 0.300 4.340 0.740 ;
        RECT  1.780 0.300 1.980 0.580 ;
        RECT  3.420 0.300 3.580 0.700 ;
        RECT  2.740 0.540 3.580 0.700 ;
        RECT  5.710 0.330 5.870 0.700 ;
        RECT  4.850 0.330 5.010 0.740 ;
        RECT  4.180 0.580 5.010 0.740 ;
        RECT  6.350 0.620 6.550 1.000 ;
        RECT  6.350 0.840 7.570 1.000 ;
        RECT  7.370 0.840 7.570 1.220 ;
        RECT  6.350 0.620 6.540 1.430 ;
        RECT  5.990 1.260 6.540 1.430 ;
        RECT  5.990 1.260 6.190 1.920 ;
        RECT  8.230 1.510 9.160 1.670 ;
        RECT  9.000 1.510 9.160 1.870 ;
        RECT  6.370 1.760 7.630 1.920 ;
        RECT  7.470 1.760 7.630 2.100 ;
        RECT  6.370 1.760 6.570 2.100 ;
        RECT  8.230 1.510 8.390 2.100 ;
        RECT  7.470 1.940 8.390 2.100 ;
        RECT  7.990 0.620 8.390 0.820 ;
        RECT  7.990 0.620 8.150 1.350 ;
        RECT  7.830 1.190 9.540 1.350 ;
        RECT  6.850 1.160 7.050 1.600 ;
        RECT  7.830 1.190 8.070 1.780 ;
        RECT  6.850 1.440 8.070 1.600 ;
        RECT  7.790 1.440 8.070 1.780 ;
        RECT  9.380 1.190 9.540 1.800 ;
        RECT  6.030 0.300 7.000 0.460 ;
        RECT  7.670 0.300 8.710 0.460 ;
        RECT  6.840 0.300 7.000 0.640 ;
        RECT  7.670 0.300 7.830 0.640 ;
        RECT  6.840 0.480 7.830 0.640 ;
        RECT  8.550 0.300 8.710 0.990 ;
        RECT  5.170 0.650 5.450 1.020 ;
        RECT  9.710 0.620 9.910 0.990 ;
        RECT  8.550 0.830 9.910 0.990 ;
        RECT  6.030 0.300 6.190 1.020 ;
        RECT  5.170 0.860 6.190 1.020 ;
        RECT  5.170 0.650 5.420 1.320 ;
        RECT  4.960 1.120 5.420 1.320 ;
        RECT  4.960 1.120 5.160 1.770 ;
        RECT  10.500 0.630 10.780 0.850 ;
        RECT  10.500 0.630 10.660 1.910 ;
        RECT  10.500 1.750 11.940 1.910 ;
        RECT  11.660 1.750 11.940 2.100 ;
        RECT  8.870 0.300 11.200 0.460 ;
        RECT  8.870 0.300 9.070 0.580 ;
        RECT  11.040 0.300 11.200 0.820 ;
        RECT  11.040 0.660 12.460 0.820 ;
        RECT  12.300 0.660 12.460 1.270 ;
        RECT  12.300 1.070 13.260 1.270 ;
        RECT  10.070 0.300 10.230 1.350 ;
        RECT  9.880 1.190 10.080 1.760 ;
        RECT  12.840 0.450 13.040 0.820 ;
        RECT  12.840 0.660 13.680 0.820 ;
        RECT  13.520 1.060 13.940 1.260 ;
        RECT  11.840 1.030 12.040 1.590 ;
        RECT  13.520 0.660 13.680 1.590 ;
        RECT  11.840 1.430 13.680 1.590 ;
        RECT  12.840 1.430 13.040 2.080 ;
        LAYER VTPH ;
        RECT  9.060 1.010 10.230 2.400 ;
        RECT  6.780 1.140 10.230 2.400 ;
        RECT  0.000 1.140 4.190 2.400 ;
        RECT  0.000 1.170 5.650 2.400 ;
        RECT  6.780 1.150 14.800 2.400 ;
        RECT  11.160 1.140 14.800 2.400 ;
        RECT  0.000 1.200 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.010 ;
        RECT  0.000 0.000 9.060 1.140 ;
        RECT  10.230 0.000 14.800 1.140 ;
        RECT  10.230 0.000 11.160 1.150 ;
        RECT  4.190 0.000 6.780 1.170 ;
        RECT  5.650 0.000 6.780 1.200 ;
    END
END SDFQSM4HM

MACRO SDFQSM2HM
    CLASS CORE ;
    FOREIGN SDFQSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.516  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.460 1.080 2.660 1.280 ;
        LAYER ME2 ;
        RECT  2.440 0.840 2.700 1.380 ;
        LAYER ME1 ;
        RECT  2.460 0.940 2.740 1.380 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 1.060 3.160 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.210 0.450 13.500 2.080 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.500 0.750 10.710 1.290 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.750 1.140 1.250 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 0.720 1.250 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.690 1.840 12.890 2.540 ;
        RECT  11.670 1.840 11.870 2.540 ;
        RECT  10.550 1.830 10.830 2.540 ;
        RECT  8.180 1.830 8.470 2.540 ;
        RECT  6.660 2.080 6.940 2.540 ;
        RECT  3.960 1.640 4.120 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.650 -0.140 12.930 0.500 ;
        RECT  11.670 -0.140 11.870 0.560 ;
        RECT  11.310 -0.140 11.510 0.560 ;
        RECT  6.820 -0.140 7.100 0.320 ;
        RECT  4.030 -0.140 4.190 0.420 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.930 1.620 1.700 ;
        RECT  0.140 1.540 1.620 1.700 ;
        RECT  0.140 0.510 0.340 1.750 ;
        RECT  2.140 0.620 2.580 0.780 ;
        RECT  2.140 0.620 2.300 1.770 ;
        RECT  2.140 1.550 2.420 1.770 ;
        RECT  3.260 0.620 3.540 0.840 ;
        RECT  3.320 0.620 3.540 1.160 ;
        RECT  3.320 1.000 4.180 1.160 ;
        RECT  3.320 0.620 3.480 1.760 ;
        RECT  3.640 1.320 4.460 1.480 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  4.300 1.320 4.460 2.100 ;
        RECT  3.640 1.320 3.800 2.100 ;
        RECT  1.620 1.940 3.800 2.100 ;
        RECT  5.100 1.640 5.300 2.100 ;
        RECT  4.300 1.940 5.300 2.100 ;
        RECT  1.780 0.300 3.860 0.460 ;
        RECT  4.370 0.330 5.390 0.490 ;
        RECT  3.700 0.300 3.860 0.740 ;
        RECT  1.780 0.300 1.980 0.650 ;
        RECT  5.230 0.330 5.390 0.700 ;
        RECT  4.370 0.330 4.530 0.740 ;
        RECT  3.700 0.580 4.530 0.740 ;
        RECT  5.870 0.620 6.070 1.000 ;
        RECT  5.870 0.840 7.160 1.000 ;
        RECT  6.960 0.840 7.160 1.220 ;
        RECT  5.870 0.620 6.060 1.430 ;
        RECT  5.620 1.260 6.060 1.430 ;
        RECT  5.620 1.260 5.820 1.920 ;
        RECT  7.860 1.510 8.790 1.670 ;
        RECT  8.630 1.510 8.790 1.870 ;
        RECT  6.000 1.760 7.260 1.920 ;
        RECT  7.100 1.760 7.260 2.100 ;
        RECT  6.000 1.760 6.200 2.100 ;
        RECT  7.860 1.510 8.020 2.100 ;
        RECT  7.100 1.940 8.020 2.100 ;
        RECT  7.620 0.620 7.980 0.820 ;
        RECT  7.620 0.620 7.780 1.350 ;
        RECT  7.420 1.190 9.170 1.350 ;
        RECT  6.480 1.160 6.680 1.600 ;
        RECT  6.480 1.440 7.700 1.600 ;
        RECT  7.420 1.190 7.700 1.780 ;
        RECT  9.010 1.190 9.170 1.800 ;
        RECT  5.550 0.300 6.630 0.460 ;
        RECT  7.260 0.300 8.300 0.460 ;
        RECT  6.470 0.300 6.630 0.640 ;
        RECT  7.260 0.300 7.420 0.640 ;
        RECT  6.470 0.480 7.420 0.640 ;
        RECT  8.140 0.300 8.300 0.990 ;
        RECT  4.690 0.650 4.970 1.020 ;
        RECT  9.300 0.620 9.500 0.990 ;
        RECT  8.140 0.830 9.500 0.990 ;
        RECT  5.550 0.300 5.710 1.020 ;
        RECT  4.690 0.860 5.710 1.020 ;
        RECT  4.690 0.650 4.930 1.400 ;
        RECT  4.620 1.120 4.820 1.780 ;
        RECT  10.060 0.620 10.340 0.840 ;
        RECT  10.130 0.620 10.340 1.610 ;
        RECT  10.130 1.450 11.150 1.610 ;
        RECT  10.130 0.620 10.290 1.780 ;
        RECT  10.990 1.450 11.150 1.990 ;
        RECT  10.990 1.830 11.390 1.990 ;
        RECT  8.460 0.300 11.130 0.460 ;
        RECT  8.460 0.300 8.660 0.580 ;
        RECT  10.970 0.300 11.130 0.880 ;
        RECT  10.970 0.720 11.870 0.880 ;
        RECT  11.710 0.720 11.870 1.180 ;
        RECT  11.710 0.980 12.110 1.180 ;
        RECT  9.660 0.300 9.820 1.350 ;
        RECT  9.510 1.190 9.710 1.760 ;
        RECT  12.210 0.450 12.410 0.820 ;
        RECT  12.210 0.660 13.050 0.820 ;
        RECT  11.310 1.040 11.510 1.500 ;
        RECT  12.890 0.660 13.050 1.500 ;
        RECT  11.310 1.340 13.050 1.500 ;
        RECT  12.210 1.340 12.410 2.080 ;
        LAYER VTPH ;
        RECT  8.650 1.080 9.810 2.400 ;
        RECT  0.000 1.140 3.710 2.400 ;
        RECT  0.000 1.170 5.170 2.400 ;
        RECT  6.410 1.140 13.600 2.400 ;
        RECT  0.000 1.200 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.080 ;
        RECT  0.000 0.000 8.650 1.140 ;
        RECT  9.810 0.000 13.600 1.140 ;
        RECT  3.710 0.000 6.410 1.170 ;
        RECT  5.170 0.000 6.410 1.200 ;
    END
END SDFQSM2HM

MACRO SDFQSM1HM
    CLASS CORE ;
    FOREIGN SDFQSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.391  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.960 1.000 2.160 1.200 ;
        LAYER ME2 ;
        RECT  1.960 0.840 2.300 1.300 ;
        LAYER ME1 ;
        RECT  1.920 0.940 2.200 1.380 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.850 1.060 3.100 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.210 0.330 13.500 2.000 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.610 0.840 11.110 1.160 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.750 1.140 1.250 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 0.720 1.250 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.690 1.840 12.890 2.540 ;
        RECT  11.670 1.840 11.870 2.540 ;
        RECT  10.550 1.830 10.830 2.540 ;
        RECT  8.180 1.830 8.470 2.540 ;
        RECT  6.660 2.080 6.940 2.540 ;
        RECT  3.960 1.640 4.120 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.650 -0.140 12.930 0.500 ;
        RECT  11.670 -0.140 11.870 0.560 ;
        RECT  6.820 -0.140 7.100 0.320 ;
        RECT  4.030 -0.140 4.190 0.420 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.930 1.620 1.700 ;
        RECT  2.460 0.820 2.620 1.700 ;
        RECT  0.140 1.540 2.620 1.700 ;
        RECT  0.140 0.530 0.340 1.750 ;
        RECT  3.260 0.620 3.540 0.840 ;
        RECT  3.320 0.620 3.540 1.160 ;
        RECT  3.320 1.000 4.180 1.160 ;
        RECT  3.320 0.620 3.480 1.760 ;
        RECT  3.640 1.320 4.460 1.480 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  4.300 1.320 4.460 2.100 ;
        RECT  3.640 1.320 3.800 2.100 ;
        RECT  1.620 1.940 3.800 2.100 ;
        RECT  5.100 1.640 5.300 2.100 ;
        RECT  4.300 1.940 5.300 2.100 ;
        RECT  1.780 0.300 3.860 0.460 ;
        RECT  4.370 0.330 5.390 0.490 ;
        RECT  3.700 0.300 3.860 0.740 ;
        RECT  1.780 0.300 1.980 0.660 ;
        RECT  5.230 0.330 5.390 0.700 ;
        RECT  4.370 0.330 4.530 0.740 ;
        RECT  3.700 0.580 4.530 0.740 ;
        RECT  5.870 0.620 6.070 1.000 ;
        RECT  5.870 0.840 7.160 1.000 ;
        RECT  6.960 0.840 7.160 1.220 ;
        RECT  5.870 0.620 6.060 1.430 ;
        RECT  5.620 1.260 6.060 1.430 ;
        RECT  5.620 1.260 5.820 1.920 ;
        RECT  7.860 1.510 8.790 1.670 ;
        RECT  8.630 1.510 8.790 1.870 ;
        RECT  6.000 1.760 7.260 1.920 ;
        RECT  7.100 1.760 7.260 2.100 ;
        RECT  6.000 1.760 6.200 2.100 ;
        RECT  7.860 1.510 8.020 2.100 ;
        RECT  7.100 1.940 8.020 2.100 ;
        RECT  7.620 0.620 7.980 0.820 ;
        RECT  7.620 0.620 7.780 1.350 ;
        RECT  7.420 1.190 9.170 1.350 ;
        RECT  6.480 1.160 6.680 1.600 ;
        RECT  6.480 1.440 7.700 1.600 ;
        RECT  7.420 1.190 7.700 1.780 ;
        RECT  9.010 1.190 9.170 1.800 ;
        RECT  5.550 0.300 6.630 0.460 ;
        RECT  7.260 0.300 8.300 0.460 ;
        RECT  6.470 0.300 6.630 0.640 ;
        RECT  7.260 0.300 7.420 0.640 ;
        RECT  6.470 0.480 7.420 0.640 ;
        RECT  8.140 0.300 8.300 0.990 ;
        RECT  4.690 0.650 4.970 1.020 ;
        RECT  9.300 0.620 9.500 0.990 ;
        RECT  8.140 0.830 9.500 0.990 ;
        RECT  5.550 0.300 5.710 1.020 ;
        RECT  4.690 0.860 5.710 1.020 ;
        RECT  4.690 0.650 4.930 1.400 ;
        RECT  4.620 1.120 4.820 1.780 ;
        RECT  10.090 0.620 10.370 1.610 ;
        RECT  10.090 1.450 11.150 1.610 ;
        RECT  10.090 0.620 10.290 1.780 ;
        RECT  10.990 1.450 11.150 1.990 ;
        RECT  10.990 1.830 11.390 1.990 ;
        RECT  8.460 0.300 11.510 0.460 ;
        RECT  8.460 0.300 8.660 0.580 ;
        RECT  11.350 0.300 11.510 0.880 ;
        RECT  11.350 0.720 11.870 0.880 ;
        RECT  11.710 0.720 11.870 1.180 ;
        RECT  11.710 0.980 12.110 1.180 ;
        RECT  9.660 0.300 9.820 1.350 ;
        RECT  9.510 1.190 9.710 1.760 ;
        RECT  12.210 0.450 12.410 0.820 ;
        RECT  12.210 0.660 13.050 0.820 ;
        RECT  11.310 1.040 11.510 1.500 ;
        RECT  12.890 0.660 13.050 1.500 ;
        RECT  11.310 1.340 13.050 1.500 ;
        RECT  12.210 1.340 12.410 2.080 ;
        LAYER VTPH ;
        RECT  1.600 1.050 2.590 2.400 ;
        RECT  8.650 1.020 9.850 2.400 ;
        RECT  0.000 1.140 3.710 2.400 ;
        RECT  0.000 1.170 5.170 2.400 ;
        RECT  6.410 1.140 13.600 2.400 ;
        RECT  0.000 1.200 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.020 ;
        RECT  0.000 0.000 8.650 1.050 ;
        RECT  0.000 0.000 1.600 1.140 ;
        RECT  2.590 0.000 8.650 1.140 ;
        RECT  9.850 0.000 13.600 1.140 ;
        RECT  3.710 0.000 6.410 1.170 ;
        RECT  5.170 0.000 6.410 1.200 ;
    END
END SDFQSM1HM

MACRO SDFQRXM2HM
    CLASS CORE ;
    FOREIGN SDFQRXM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.417  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.170 1.050 1.370 1.250 ;
        LAYER ME2 ;
        RECT  1.170 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.000 0.970 1.470 1.300 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.740 1.300 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.468  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.820 2.950 7.100 4.360 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.840 4.100 5.280 4.480 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.670 3.670 1.160 3.900 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 3.440 2.580 3.720 ;
        RECT  1.700 3.440 1.900 3.960 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.280 2.260 6.480 3.270 ;
        RECT  4.830 1.760 5.110 2.540 ;
        RECT  4.420 2.260 4.700 2.770 ;
        RECT  0.660 2.200 0.940 2.540 ;
        RECT  0.620 2.260 0.900 3.160 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.880 -0.140 7.100 0.870 ;
        RECT  4.870 -0.140 5.070 0.610 ;
        RECT  0.680 -0.140 0.880 0.390 ;
        RECT  0.000 4.660 7.200 4.940 ;
        RECT  6.260 4.480 6.540 4.940 ;
        RECT  5.440 3.960 5.600 4.940 ;
        RECT  0.620 4.060 0.900 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.320 1.540 3.480 ;
        RECT  1.380 3.320 1.540 3.930 ;
        RECT  0.140 2.940 0.340 4.270 ;
        RECT  0.920 0.650 1.790 0.810 ;
        RECT  1.630 1.020 1.930 1.220 ;
        RECT  1.630 0.650 1.790 1.720 ;
        RECT  0.920 1.560 1.790 1.720 ;
        RECT  0.140 0.390 0.340 2.040 ;
        RECT  0.140 1.880 2.720 2.040 ;
        RECT  2.420 1.880 2.720 2.100 ;
        RECT  2.030 3.120 2.900 3.280 ;
        RECT  2.740 3.120 2.900 4.040 ;
        RECT  2.260 3.880 2.900 4.040 ;
        RECT  2.260 3.880 2.540 4.160 ;
        RECT  1.580 2.720 2.900 2.880 ;
        RECT  2.620 2.720 2.900 2.960 ;
        RECT  1.580 2.720 1.780 3.100 ;
        RECT  1.740 4.200 1.940 4.480 ;
        RECT  2.780 4.200 2.980 4.480 ;
        RECT  1.740 4.320 2.980 4.480 ;
        RECT  1.990 0.600 2.310 0.800 ;
        RECT  2.140 0.600 2.310 1.660 ;
        RECT  2.030 1.440 2.310 1.660 ;
        RECT  2.030 1.500 3.060 1.660 ;
        RECT  2.900 1.500 3.060 2.070 ;
        RECT  2.900 1.910 4.360 2.070 ;
        RECT  3.060 3.390 3.340 3.590 ;
        RECT  3.180 3.390 3.340 4.480 ;
        RECT  3.180 4.320 4.520 4.480 ;
        RECT  2.510 0.320 4.710 0.480 ;
        RECT  2.510 0.320 2.710 1.220 ;
        RECT  2.510 1.060 3.420 1.220 ;
        RECT  3.220 1.060 3.420 1.740 ;
        RECT  3.860 2.760 4.060 3.120 ;
        RECT  5.220 2.880 5.500 3.120 ;
        RECT  3.860 2.960 5.500 3.120 ;
        RECT  3.180 2.880 3.660 3.040 ;
        RECT  3.500 2.880 3.660 3.800 ;
        RECT  3.500 3.600 5.600 3.800 ;
        RECT  3.820 3.600 4.100 4.160 ;
        RECT  3.100 0.640 3.740 0.800 ;
        RECT  3.580 0.640 3.740 1.280 ;
        RECT  3.580 1.120 5.810 1.280 ;
        RECT  3.740 1.120 3.940 1.740 ;
        RECT  5.740 2.990 5.940 3.440 ;
        RECT  4.160 3.280 5.940 3.440 ;
        RECT  5.780 2.990 5.940 4.200 ;
        RECT  5.780 4.000 6.180 4.200 ;
        RECT  3.940 0.640 4.220 0.960 ;
        RECT  6.200 0.680 6.500 0.960 ;
        RECT  3.940 0.800 6.500 0.960 ;
        RECT  4.260 1.440 6.640 1.600 ;
        RECT  6.360 1.440 6.640 1.720 ;
        RECT  4.260 1.440 4.460 1.750 ;
        RECT  5.630 0.300 6.640 0.500 ;
        RECT  5.350 1.760 5.630 2.100 ;
        RECT  5.350 1.940 6.650 2.100 ;
        LAYER VTPH ;
        RECT  1.790 1.140 2.630 3.640 ;
        RECT  0.000 1.140 0.850 3.660 ;
        RECT  1.790 1.160 5.890 3.640 ;
        RECT  4.470 1.090 5.890 3.640 ;
        RECT  0.000 1.200 7.200 3.640 ;
        RECT  0.000 1.190 1.900 3.660 ;
        RECT  6.350 1.200 7.200 3.660 ;
        LAYER VTNH ;
        RECT  1.900 3.640 6.350 4.800 ;
        RECT  0.000 3.660 7.200 4.800 ;
        RECT  0.000 0.000 7.200 1.090 ;
        RECT  0.000 0.000 4.470 1.140 ;
        RECT  2.630 0.000 4.470 1.160 ;
        RECT  0.850 0.000 1.790 1.190 ;
        RECT  5.890 0.000 7.200 1.200 ;
    END
END SDFQRXM2HM

MACRO SDFQRSM8HM
    CLASS CORE ;
    FOREIGN SDFQRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.497  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.190 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.968  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.400 0.850 17.600 2.080 ;
        RECT  17.420 0.410 17.600 2.080 ;
        RECT  16.360 0.850 17.600 1.100 ;
        RECT  16.360 0.450 16.560 2.080 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.319  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.226  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 10.280  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.980 0.800 13.260 1.060 ;
        RECT  12.000 0.800 13.260 0.960 ;
        RECT  12.000 0.800 12.300 1.240 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.990 0.900 15.560 1.160 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.061  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.400 2.540 ;
        RECT  17.920 1.480 18.120 2.540 ;
        RECT  16.880 1.840 17.080 2.540 ;
        RECT  15.780 2.020 15.980 2.540 ;
        RECT  14.540 1.860 14.820 2.540 ;
        RECT  13.400 1.860 13.680 2.540 ;
        RECT  12.320 1.800 12.520 2.540 ;
        RECT  8.920 2.080 9.200 2.540 ;
        RECT  4.360 1.980 4.520 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.400 0.140 ;
        RECT  17.920 -0.140 18.120 0.730 ;
        RECT  16.880 -0.140 17.080 0.560 ;
        RECT  15.740 -0.140 16.020 0.320 ;
        RECT  14.340 -0.140 14.620 0.320 ;
        RECT  12.220 -0.140 12.500 0.320 ;
        RECT  7.900 -0.140 8.100 0.400 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.770 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.260 ;
        RECT  3.700 1.100 4.860 1.260 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.660 4.840 1.820 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.680 1.660 4.840 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.660 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.680 1.940 5.660 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.620 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.620 5.460 1.510 ;
        RECT  5.000 1.350 5.460 1.510 ;
        RECT  5.000 1.350 5.160 1.780 ;
        RECT  6.720 1.620 8.160 1.780 ;
        RECT  6.460 0.900 8.800 1.060 ;
        RECT  8.640 0.900 8.800 1.260 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  5.980 1.240 6.660 1.400 ;
        RECT  5.980 1.240 6.180 2.020 ;
        RECT  8.960 0.620 9.700 0.780 ;
        RECT  6.930 1.240 8.480 1.400 ;
        RECT  8.320 1.240 8.480 1.600 ;
        RECT  8.960 0.620 9.120 1.600 ;
        RECT  8.320 1.440 9.880 1.600 ;
        RECT  9.680 1.440 9.880 1.760 ;
        RECT  8.320 1.760 9.520 1.920 ;
        RECT  9.360 1.760 9.520 2.100 ;
        RECT  8.320 1.760 8.480 2.100 ;
        RECT  6.340 1.940 8.480 2.100 ;
        RECT  10.080 1.660 10.240 2.100 ;
        RECT  9.360 1.940 10.240 2.100 ;
        RECT  9.720 1.080 11.200 1.280 ;
        RECT  8.260 0.300 11.240 0.460 ;
        RECT  7.460 0.300 7.740 0.720 ;
        RECT  8.260 0.300 8.420 0.720 ;
        RECT  7.460 0.560 8.420 0.720 ;
        RECT  9.980 0.620 10.260 0.900 ;
        RECT  9.980 0.740 11.520 0.900 ;
        RECT  12.460 1.120 12.780 1.380 ;
        RECT  14.120 1.120 14.400 1.380 ;
        RECT  12.460 1.220 14.400 1.380 ;
        RECT  12.460 1.120 12.620 1.640 ;
        RECT  12.000 1.480 12.620 1.640 ;
        RECT  10.780 1.510 11.520 1.710 ;
        RECT  11.360 0.740 11.520 2.100 ;
        RECT  11.350 1.510 11.520 2.100 ;
        RECT  12.000 1.480 12.160 2.100 ;
        RECT  11.350 1.940 12.160 2.100 ;
        RECT  13.420 0.620 13.700 0.960 ;
        RECT  13.420 0.800 14.720 0.960 ;
        RECT  15.720 0.980 15.880 1.480 ;
        RECT  14.560 1.320 15.880 1.480 ;
        RECT  14.560 0.800 14.720 1.700 ;
        RECT  12.800 1.540 14.720 1.700 ;
        RECT  12.660 0.300 14.100 0.460 ;
        RECT  13.940 0.300 14.100 0.640 ;
        RECT  14.820 0.400 15.100 0.640 ;
        RECT  12.660 0.300 12.820 0.640 ;
        RECT  11.680 0.480 12.820 0.640 ;
        RECT  13.940 0.480 16.200 0.640 ;
        RECT  11.680 0.480 11.840 1.780 ;
        RECT  16.040 0.480 16.200 1.860 ;
        RECT  15.100 1.700 16.200 1.860 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  9.820 1.080 10.020 1.280 ;
        LAYER ME2 ;
        RECT  6.720 0.400 10.020 0.600 ;
        RECT  9.820 0.400 10.020 1.380 ;
        LAYER VTPH ;
        RECT  7.070 1.080 9.200 2.400 ;
        RECT  12.220 1.080 13.070 2.400 ;
        RECT  0.000 1.140 5.660 2.400 ;
        RECT  7.070 1.140 18.400 2.400 ;
        RECT  0.000 1.200 18.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.400 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.200 0.000 12.220 1.140 ;
        RECT  13.070 0.000 18.400 1.140 ;
        RECT  5.660 0.000 7.070 1.200 ;
    END
END SDFQRSM8HM

MACRO SDFQRSM4HM
    CLASS CORE ;
    FOREIGN SDFQRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 16.075  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.940 0.400 11.140 0.600 ;
        LAYER ME2 ;
        RECT  10.800 0.400 11.240 0.760 ;
        LAYER ME1 ;
        RECT  10.800 0.300 11.240 0.600 ;
        RECT  8.260 0.300 11.240 0.460 ;
        RECT  7.460 0.560 8.420 0.720 ;
        RECT  8.260 0.300 8.420 0.720 ;
        RECT  7.460 0.300 7.740 0.720 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.521  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.160 0.780 15.500 1.280 ;
        RECT  15.160 0.410 15.360 2.080 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.910 0.900 14.360 1.160 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.000 2.540 ;
        RECT  15.660 1.480 15.860 2.540 ;
        RECT  14.520 2.080 14.800 2.540 ;
        RECT  13.460 1.860 13.740 2.540 ;
        RECT  12.380 1.580 12.660 2.540 ;
        RECT  8.920 2.080 9.200 2.540 ;
        RECT  4.360 1.980 4.520 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.000 0.140 ;
        RECT  15.660 -0.140 15.860 0.730 ;
        RECT  14.510 -0.140 14.790 0.320 ;
        RECT  13.260 -0.140 13.540 0.320 ;
        RECT  7.900 -0.140 8.100 0.400 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.300 ;
        RECT  3.700 1.100 4.820 1.300 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.660 4.840 1.820 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.680 1.660 4.840 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.660 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.680 1.940 5.660 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.640 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.640 5.460 1.510 ;
        RECT  5.000 1.350 5.460 1.510 ;
        RECT  5.000 1.350 5.160 1.780 ;
        RECT  6.720 1.620 8.160 1.780 ;
        RECT  6.460 0.900 8.800 1.060 ;
        RECT  8.640 0.900 8.800 1.260 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  5.980 1.240 6.660 1.400 ;
        RECT  5.980 1.240 6.180 2.020 ;
        RECT  8.960 0.620 9.700 0.780 ;
        RECT  6.930 1.240 8.480 1.400 ;
        RECT  8.320 1.240 8.480 1.600 ;
        RECT  8.960 0.620 9.120 1.600 ;
        RECT  8.320 1.440 9.880 1.600 ;
        RECT  9.680 1.440 9.880 1.760 ;
        RECT  8.320 1.760 9.520 1.920 ;
        RECT  9.360 1.760 9.520 2.100 ;
        RECT  8.320 1.760 8.480 2.100 ;
        RECT  6.340 1.940 8.480 2.100 ;
        RECT  10.080 1.660 10.240 2.100 ;
        RECT  9.360 1.940 10.240 2.100 ;
        RECT  9.720 1.080 11.200 1.280 ;
        RECT  10.020 0.620 10.300 0.920 ;
        RECT  10.020 0.760 11.520 0.920 ;
        RECT  13.040 1.120 13.320 1.380 ;
        RECT  12.000 1.220 13.320 1.380 ;
        RECT  10.780 1.510 11.520 1.710 ;
        RECT  11.360 0.760 11.520 2.100 ;
        RECT  11.350 1.510 11.520 2.100 ;
        RECT  12.000 1.220 12.160 2.100 ;
        RECT  11.350 1.940 12.160 2.100 ;
        RECT  12.380 0.620 12.660 0.960 ;
        RECT  12.380 0.800 13.640 0.960 ;
        RECT  14.520 0.980 14.680 1.480 ;
        RECT  13.480 1.320 14.680 1.480 ;
        RECT  13.480 0.800 13.640 1.700 ;
        RECT  12.860 1.540 13.640 1.700 ;
        RECT  11.680 0.300 13.020 0.460 ;
        RECT  12.860 0.300 13.020 0.640 ;
        RECT  12.860 0.480 15.000 0.640 ;
        RECT  11.680 0.300 11.840 1.780 ;
        RECT  14.840 0.480 15.000 1.800 ;
        RECT  14.020 1.640 15.000 1.800 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  9.820 1.080 10.020 1.280 ;
        LAYER ME2 ;
        RECT  6.720 0.400 10.020 0.600 ;
        RECT  9.820 0.400 10.020 1.380 ;
        LAYER VTPH ;
        RECT  7.070 1.080 9.200 2.400 ;
        RECT  0.000 1.140 4.090 2.400 ;
        RECT  0.000 1.160 5.660 2.400 ;
        RECT  7.070 1.140 16.000 2.400 ;
        RECT  0.000 1.200 16.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.000 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.200 0.000 16.000 1.140 ;
        RECT  4.090 0.000 7.070 1.160 ;
        RECT  5.660 0.000 7.070 1.200 ;
    END
END SDFQRSM4HM

MACRO SDFQRSM2HM
    CLASS CORE ;
    FOREIGN SDFQRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.600 1.060 2.800 1.260 ;
        LAYER ME2 ;
        RECT  2.440 0.900 2.860 1.280 ;
        LAYER ME1 ;
        RECT  2.540 1.040 2.860 1.400 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 16.075  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.940 0.400 11.140 0.600 ;
        LAYER ME2 ;
        RECT  10.800 0.400 11.240 0.760 ;
        LAYER ME1 ;
        RECT  10.800 0.300 11.240 0.600 ;
        RECT  8.260 0.300 11.240 0.460 ;
        RECT  7.460 0.560 8.420 0.720 ;
        RECT  8.260 0.300 8.420 0.720 ;
        RECT  7.460 0.300 7.740 0.720 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.040 3.500 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.160 0.780 15.500 1.280 ;
        RECT  15.160 0.410 15.360 2.080 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.910 0.900 14.360 1.160 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.850 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  14.520 2.080 14.800 2.540 ;
        RECT  13.460 1.860 13.740 2.540 ;
        RECT  12.380 1.580 12.660 2.540 ;
        RECT  8.920 2.080 9.200 2.540 ;
        RECT  4.360 1.980 4.520 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  14.510 -0.140 14.790 0.320 ;
        RECT  13.260 -0.140 13.540 0.320 ;
        RECT  7.900 -0.140 8.100 0.400 ;
        RECT  4.580 -0.140 4.780 0.600 ;
        RECT  3.140 -0.140 3.340 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.050 1.640 1.640 ;
        RECT  0.140 1.480 1.640 1.640 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  2.160 0.620 2.660 0.780 ;
        RECT  2.160 0.620 2.320 1.780 ;
        RECT  2.160 1.580 2.440 1.780 ;
        RECT  3.820 0.620 4.100 1.300 ;
        RECT  3.700 1.100 4.820 1.300 ;
        RECT  3.700 1.100 3.860 1.760 ;
        RECT  4.020 1.660 4.840 1.820 ;
        RECT  2.600 1.760 3.540 1.920 ;
        RECT  1.620 1.860 1.900 2.100 ;
        RECT  3.380 1.760 3.540 2.100 ;
        RECT  4.680 1.660 4.840 2.100 ;
        RECT  2.600 1.760 2.760 2.100 ;
        RECT  1.620 1.940 2.760 2.100 ;
        RECT  4.020 1.660 4.200 2.100 ;
        RECT  3.380 1.940 4.200 2.100 ;
        RECT  5.460 1.740 5.660 2.100 ;
        RECT  4.680 1.940 5.660 2.100 ;
        RECT  1.840 0.300 2.980 0.460 ;
        RECT  3.500 0.300 4.420 0.460 ;
        RECT  4.940 0.300 5.980 0.460 ;
        RECT  5.780 0.300 5.980 0.600 ;
        RECT  2.820 0.300 2.980 0.880 ;
        RECT  1.840 0.300 2.000 0.740 ;
        RECT  4.260 0.300 4.420 0.920 ;
        RECT  3.500 0.300 3.660 0.880 ;
        RECT  2.820 0.720 3.660 0.880 ;
        RECT  4.940 0.300 5.100 0.920 ;
        RECT  4.260 0.760 5.100 0.920 ;
        RECT  6.140 0.300 7.020 0.460 ;
        RECT  6.820 0.300 7.020 0.720 ;
        RECT  5.260 0.640 5.540 0.920 ;
        RECT  6.140 0.300 6.300 0.920 ;
        RECT  5.260 0.760 6.300 0.920 ;
        RECT  5.260 0.640 5.460 1.510 ;
        RECT  5.000 1.350 5.460 1.510 ;
        RECT  5.000 1.350 5.160 1.780 ;
        RECT  6.720 1.620 8.160 1.780 ;
        RECT  6.460 0.900 8.800 1.060 ;
        RECT  8.640 0.900 8.800 1.260 ;
        RECT  6.460 0.620 6.660 1.400 ;
        RECT  5.980 1.240 6.660 1.400 ;
        RECT  5.980 1.240 6.180 2.020 ;
        RECT  8.960 0.620 9.700 0.780 ;
        RECT  6.930 1.240 8.480 1.400 ;
        RECT  8.320 1.240 8.480 1.600 ;
        RECT  8.960 0.620 9.120 1.600 ;
        RECT  8.320 1.440 9.880 1.600 ;
        RECT  9.680 1.440 9.880 1.760 ;
        RECT  8.320 1.760 9.520 1.920 ;
        RECT  9.360 1.760 9.520 2.100 ;
        RECT  8.320 1.760 8.480 2.100 ;
        RECT  6.340 1.940 8.480 2.100 ;
        RECT  10.080 1.660 10.240 2.100 ;
        RECT  9.360 1.940 10.240 2.100 ;
        RECT  9.720 1.080 11.200 1.280 ;
        RECT  10.020 0.620 10.300 0.920 ;
        RECT  10.020 0.760 11.520 0.920 ;
        RECT  13.040 1.120 13.320 1.380 ;
        RECT  12.000 1.220 13.320 1.380 ;
        RECT  10.780 1.510 11.520 1.710 ;
        RECT  11.360 0.760 11.520 2.100 ;
        RECT  11.350 1.510 11.520 2.100 ;
        RECT  12.000 1.220 12.160 2.100 ;
        RECT  11.350 1.940 12.160 2.100 ;
        RECT  12.380 0.620 12.660 0.960 ;
        RECT  12.380 0.800 13.640 0.960 ;
        RECT  14.520 0.980 14.680 1.480 ;
        RECT  13.480 1.320 14.680 1.480 ;
        RECT  13.480 0.800 13.640 1.700 ;
        RECT  12.860 1.540 13.640 1.700 ;
        RECT  11.680 0.300 13.020 0.460 ;
        RECT  12.860 0.300 13.020 0.640 ;
        RECT  12.860 0.480 15.000 0.640 ;
        RECT  11.680 0.300 11.840 1.780 ;
        RECT  14.840 0.480 15.000 1.800 ;
        RECT  14.020 1.640 15.000 1.800 ;
        LAYER VI1 ;
        RECT  6.820 0.400 7.020 0.600 ;
        RECT  9.820 1.080 10.020 1.280 ;
        LAYER ME2 ;
        RECT  6.720 0.400 10.020 0.600 ;
        RECT  9.820 0.400 10.020 1.380 ;
        LAYER VTPH ;
        RECT  7.070 1.080 9.200 2.400 ;
        RECT  0.000 1.140 4.090 2.400 ;
        RECT  0.000 1.160 5.660 2.400 ;
        RECT  7.070 1.140 15.600 2.400 ;
        RECT  0.000 1.200 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.080 ;
        RECT  0.000 0.000 7.070 1.140 ;
        RECT  9.200 0.000 15.600 1.140 ;
        RECT  4.090 0.000 7.070 1.160 ;
        RECT  5.660 0.000 7.070 1.200 ;
    END
END SDFQRSM2HM

MACRO SDFQRSM1HM
    CLASS CORE ;
    FOREIGN SDFQRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.345  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 15.761  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 21.772  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  12.550 0.950 12.750 1.150 ;
        LAYER ME2 ;
        RECT  12.500 0.840 12.770 1.350 ;
        LAYER ME1 ;
        RECT  12.520 0.800 12.780 1.260 ;
        RECT  11.580 0.800 12.780 0.960 ;
        RECT  11.580 0.800 11.860 1.020 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.344  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.930 0.960 2.130 1.160 ;
        LAYER ME2 ;
        RECT  1.930 0.840 2.300 1.280 ;
        LAYER ME1 ;
        RECT  1.800 0.900 2.190 1.220 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.840 3.160 1.300 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.860 0.440 15.100 1.860 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.540 1.160 13.960 1.500 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.260 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.480 1.640 0.870 ;
        RECT  0.500 0.480 1.640 0.640 ;
        RECT  0.500 0.480 0.700 1.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.260 2.020 14.460 2.540 ;
        RECT  12.980 1.860 13.260 2.540 ;
        RECT  11.900 1.520 12.100 2.540 ;
        RECT  8.550 2.080 8.830 2.540 ;
        RECT  4.150 2.020 4.350 2.540 ;
        RECT  2.680 2.020 2.880 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.240 -0.140 14.520 0.320 ;
        RECT  11.860 -0.140 12.140 0.320 ;
        RECT  7.530 -0.140 7.810 0.420 ;
        RECT  4.130 -0.140 4.330 0.600 ;
        RECT  2.660 -0.140 2.940 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.440 1.380 2.680 1.540 ;
        RECT  2.480 0.850 2.680 1.540 ;
        RECT  1.440 1.070 1.640 1.700 ;
        RECT  0.140 1.540 1.640 1.700 ;
        RECT  0.140 0.300 0.340 1.820 ;
        RECT  3.420 1.100 4.610 1.300 ;
        RECT  3.420 0.620 3.620 1.780 ;
        RECT  1.950 1.700 3.200 1.860 ;
        RECT  3.810 1.700 4.670 1.860 ;
        RECT  3.040 1.700 3.200 2.100 ;
        RECT  4.510 1.700 4.670 2.100 ;
        RECT  1.580 1.860 2.110 2.020 ;
        RECT  3.810 1.700 3.990 2.100 ;
        RECT  3.040 1.940 3.990 2.100 ;
        RECT  5.310 1.740 5.510 2.100 ;
        RECT  4.510 1.940 5.510 2.100 ;
        RECT  3.100 0.300 3.970 0.460 ;
        RECT  4.490 0.300 5.550 0.460 ;
        RECT  1.820 0.370 2.020 0.680 ;
        RECT  5.350 0.300 5.550 0.600 ;
        RECT  3.100 0.300 3.260 0.680 ;
        RECT  1.820 0.520 3.260 0.680 ;
        RECT  3.810 0.300 3.970 0.920 ;
        RECT  4.490 0.300 4.650 0.920 ;
        RECT  3.810 0.760 4.650 0.920 ;
        RECT  5.710 0.300 6.670 0.460 ;
        RECT  6.470 0.300 6.670 0.720 ;
        RECT  4.830 0.640 5.110 0.920 ;
        RECT  5.710 0.300 5.870 0.920 ;
        RECT  4.830 0.760 5.870 0.920 ;
        RECT  4.830 0.640 5.030 1.780 ;
        RECT  6.390 1.560 7.750 1.780 ;
        RECT  6.030 0.920 7.950 1.080 ;
        RECT  6.030 0.680 6.310 1.400 ;
        RECT  5.830 1.240 6.030 2.020 ;
        RECT  8.630 0.620 9.330 0.780 ;
        RECT  6.710 1.240 8.110 1.400 ;
        RECT  7.950 1.240 8.110 1.600 ;
        RECT  8.630 0.620 8.790 1.600 ;
        RECT  7.950 1.440 9.520 1.600 ;
        RECT  9.320 1.440 9.520 1.780 ;
        RECT  7.950 1.760 9.160 1.920 ;
        RECT  9.000 1.760 9.160 2.100 ;
        RECT  7.950 1.760 8.110 2.100 ;
        RECT  6.190 1.940 8.110 2.100 ;
        RECT  9.720 1.660 9.880 2.100 ;
        RECT  9.000 1.940 9.880 2.100 ;
        RECT  10.580 1.000 10.780 1.280 ;
        RECT  9.350 1.080 10.780 1.280 ;
        RECT  7.970 0.300 10.880 0.460 ;
        RECT  7.090 0.300 7.370 0.740 ;
        RECT  7.970 0.300 8.130 0.740 ;
        RECT  7.090 0.580 8.130 0.740 ;
        RECT  9.710 0.620 9.990 0.820 ;
        RECT  9.710 0.660 11.100 0.820 ;
        RECT  12.080 1.120 12.360 1.340 ;
        RECT  11.580 1.180 12.360 1.340 ;
        RECT  10.420 1.500 11.100 1.700 ;
        RECT  10.940 0.660 11.100 2.100 ;
        RECT  10.930 1.500 11.100 2.100 ;
        RECT  11.580 1.180 11.740 2.100 ;
        RECT  10.930 1.940 11.740 2.100 ;
        RECT  12.940 0.620 13.220 0.960 ;
        RECT  12.940 0.800 14.360 0.960 ;
        RECT  14.160 0.800 14.360 1.300 ;
        RECT  12.940 0.620 13.100 1.700 ;
        RECT  12.420 1.500 13.100 1.700 ;
        RECT  12.300 0.300 13.660 0.460 ;
        RECT  13.460 0.300 13.660 0.640 ;
        RECT  12.300 0.300 12.460 0.640 ;
        RECT  11.260 0.480 12.460 0.640 ;
        RECT  13.460 0.480 14.680 0.640 ;
        RECT  11.260 0.480 11.420 1.780 ;
        RECT  14.520 0.480 14.680 1.860 ;
        RECT  13.540 1.700 14.680 1.860 ;
        LAYER VI1 ;
        RECT  6.470 0.400 6.670 0.600 ;
        RECT  9.450 1.080 9.650 1.280 ;
        LAYER ME2 ;
        RECT  6.370 0.400 9.650 0.600 ;
        RECT  9.450 0.400 9.650 1.380 ;
        LAYER VTPH ;
        RECT  7.480 1.080 8.830 2.400 ;
        RECT  1.370 1.050 2.650 2.400 ;
        RECT  0.000 1.140 2.650 2.400 ;
        RECT  7.480 1.140 15.200 2.400 ;
        RECT  0.000 1.200 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 1.050 ;
        RECT  2.650 0.000 15.200 1.080 ;
        RECT  0.000 0.000 1.370 1.140 ;
        RECT  8.830 0.000 15.200 1.140 ;
        RECT  2.650 0.000 7.480 1.200 ;
    END
END SDFQRSM1HM

MACRO SDFQRM8HM
    CLASS CORE ;
    FOREIGN SDFQRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.140 1.300 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.740 1.300 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.049  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.940 3.120 8.180 4.360 ;
        RECT  6.810 3.550 8.180 4.050 ;
        RECT  7.890 3.120 8.180 4.050 ;
        RECT  6.810 3.550 7.100 4.360 ;
        RECT  6.810 3.120 7.090 4.360 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.800 4.100 5.240 4.480 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.650 3.670 1.160 3.900 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 3.440 2.580 3.720 ;
        RECT  1.700 3.440 1.900 3.960 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.460 1.480 8.660 3.160 ;
        RECT  8.450 1.480 8.660 2.540 ;
        RECT  7.410 2.260 7.610 2.960 ;
        RECT  6.220 2.260 6.420 3.270 ;
        RECT  6.090 2.080 6.370 2.540 ;
        RECT  5.010 1.760 5.290 2.540 ;
        RECT  4.380 2.260 4.660 2.770 ;
        RECT  1.560 2.140 1.840 2.540 ;
        RECT  0.660 2.140 0.940 2.540 ;
        RECT  0.620 2.260 0.900 3.160 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.450 -0.140 8.650 0.840 ;
        RECT  6.730 -0.140 7.010 0.320 ;
        RECT  5.050 -0.140 5.250 0.610 ;
        RECT  1.660 -0.140 1.860 0.600 ;
        RECT  0.660 -0.140 0.860 0.560 ;
        RECT  0.000 4.660 8.800 4.940 ;
        RECT  8.460 4.140 8.660 4.940 ;
        RECT  7.420 4.210 7.620 4.940 ;
        RECT  6.380 4.100 6.580 4.940 ;
        RECT  5.400 4.140 5.560 4.940 ;
        RECT  0.620 4.060 0.900 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.320 1.540 3.480 ;
        RECT  1.380 3.320 1.540 3.930 ;
        RECT  0.140 2.940 0.340 4.270 ;
        RECT  1.060 0.400 1.480 0.560 ;
        RECT  1.300 0.400 1.480 1.220 ;
        RECT  1.300 1.020 2.040 1.220 ;
        RECT  1.320 0.400 1.480 1.660 ;
        RECT  0.960 1.500 1.480 1.660 ;
        RECT  0.140 0.390 0.340 1.980 ;
        RECT  0.140 1.820 2.240 1.980 ;
        RECT  2.080 1.940 2.840 2.100 ;
        RECT  2.030 3.120 2.900 3.280 ;
        RECT  2.740 3.120 2.900 4.040 ;
        RECT  2.260 3.880 2.900 4.040 ;
        RECT  2.260 3.880 2.540 4.160 ;
        RECT  1.580 2.720 2.900 2.880 ;
        RECT  2.620 2.720 2.900 2.960 ;
        RECT  1.580 2.720 1.780 3.100 ;
        RECT  1.740 4.200 1.940 4.480 ;
        RECT  2.780 4.200 2.980 4.480 ;
        RECT  1.740 4.320 2.980 4.480 ;
        RECT  3.060 3.390 3.340 3.590 ;
        RECT  3.180 3.390 3.340 4.480 ;
        RECT  3.180 4.320 4.480 4.480 ;
        RECT  2.140 0.380 2.380 0.700 ;
        RECT  2.200 0.380 2.380 1.660 ;
        RECT  2.080 1.500 3.160 1.660 ;
        RECT  3.000 1.500 3.160 2.070 ;
        RECT  3.000 1.910 4.510 2.070 ;
        RECT  2.690 0.320 4.890 0.480 ;
        RECT  2.690 0.320 2.890 1.220 ;
        RECT  2.690 1.060 3.530 1.220 ;
        RECT  3.330 1.060 3.530 1.750 ;
        RECT  3.820 2.760 4.020 3.120 ;
        RECT  5.180 2.880 5.460 3.120 ;
        RECT  3.820 2.960 5.460 3.120 ;
        RECT  3.120 2.880 3.660 3.040 ;
        RECT  3.500 2.880 3.660 3.850 ;
        RECT  3.500 3.650 5.560 3.850 ;
        RECT  3.780 3.650 4.060 4.160 ;
        RECT  5.700 2.990 5.900 3.440 ;
        RECT  4.120 3.280 5.900 3.440 ;
        RECT  5.740 2.990 5.900 4.420 ;
        RECT  5.740 4.220 6.140 4.420 ;
        RECT  3.210 0.640 3.850 0.800 ;
        RECT  3.690 0.640 3.850 1.280 ;
        RECT  3.690 1.120 6.350 1.280 ;
        RECT  3.850 1.120 4.050 1.750 ;
        RECT  4.010 0.640 4.370 0.800 ;
        RECT  7.490 0.620 7.770 0.960 ;
        RECT  4.210 0.800 7.770 0.960 ;
        RECT  4.450 1.440 7.840 1.600 ;
        RECT  7.560 1.440 7.840 1.660 ;
        RECT  4.450 1.440 4.650 1.750 ;
        RECT  7.170 0.300 8.200 0.460 ;
        RECT  7.170 0.300 7.330 0.640 ;
        RECT  5.810 0.480 7.330 0.640 ;
        RECT  5.490 1.760 7.190 1.920 ;
        RECT  8.000 0.300 8.200 1.980 ;
        RECT  7.040 1.820 8.200 1.980 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.540 3.640 ;
        RECT  4.450 1.140 8.800 3.640 ;
        RECT  0.000 1.170 8.800 3.640 ;
        RECT  0.000 1.140 1.900 3.660 ;
        RECT  4.840 1.140 8.800 3.660 ;
        LAYER VTNH ;
        RECT  1.900 3.640 4.840 4.800 ;
        RECT  0.000 3.660 8.800 4.800 ;
        RECT  0.000 0.000 8.800 1.140 ;
        RECT  2.540 0.000 4.450 1.170 ;
    END
END SDFQRM8HM

MACRO SDFQRM4HM
    CLASS CORE ;
    FOREIGN SDFQRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        ANTENNAGATEAREA 0.074  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.591  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.170 1.050 1.370 1.250 ;
        LAYER ME2 ;
        RECT  1.170 0.840 1.530 1.560 ;
        LAYER ME1 ;
        RECT  1.000 0.970 1.470 1.300 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.740 1.300 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.785  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.890 2.730 8.170 4.360 ;
        RECT  6.730 3.640 8.170 3.900 ;
        RECT  6.730 3.120 7.010 4.360 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.840 4.100 5.280 4.480 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.650 3.670 1.160 3.900 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 3.440 2.580 3.720 ;
        RECT  1.700 3.440 1.900 3.960 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  8.080 1.440 8.260 2.540 ;
        RECT  7.250 2.260 7.530 3.120 ;
        RECT  6.260 2.260 6.460 3.270 ;
        RECT  5.980 2.080 6.260 2.540 ;
        RECT  4.900 1.760 5.180 2.540 ;
        RECT  4.420 2.260 4.700 2.770 ;
        RECT  0.660 2.200 0.940 2.540 ;
        RECT  0.620 2.260 0.900 3.160 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  8.080 -0.140 8.280 0.870 ;
        RECT  6.620 -0.140 6.900 0.320 ;
        RECT  4.940 -0.140 5.140 0.610 ;
        RECT  0.680 -0.140 0.880 0.390 ;
        RECT  0.000 4.660 8.400 4.940 ;
        RECT  7.290 4.210 7.490 4.940 ;
        RECT  5.440 4.140 5.600 4.940 ;
        RECT  0.620 4.060 0.900 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.320 1.540 3.480 ;
        RECT  1.380 3.320 1.540 3.930 ;
        RECT  0.140 2.940 0.340 4.270 ;
        RECT  0.920 0.650 1.790 0.810 ;
        RECT  1.630 1.020 1.930 1.220 ;
        RECT  1.630 0.650 1.790 1.720 ;
        RECT  0.920 1.560 1.790 1.720 ;
        RECT  0.140 0.390 0.340 2.040 ;
        RECT  0.140 1.880 2.720 2.040 ;
        RECT  2.420 1.880 2.720 2.100 ;
        RECT  2.030 3.120 2.900 3.280 ;
        RECT  2.740 3.120 2.900 4.040 ;
        RECT  2.260 3.880 2.900 4.040 ;
        RECT  2.260 3.880 2.540 4.160 ;
        RECT  1.580 2.720 2.900 2.880 ;
        RECT  2.620 2.720 2.900 2.960 ;
        RECT  1.580 2.720 1.780 3.100 ;
        RECT  1.740 4.200 1.940 4.480 ;
        RECT  2.780 4.200 2.980 4.480 ;
        RECT  1.740 4.320 2.980 4.480 ;
        RECT  1.990 0.600 2.310 0.800 ;
        RECT  2.140 0.600 2.310 1.660 ;
        RECT  2.030 1.440 2.310 1.660 ;
        RECT  2.030 1.500 3.060 1.660 ;
        RECT  2.900 1.500 3.060 2.070 ;
        RECT  2.900 1.910 4.400 2.070 ;
        RECT  3.060 3.390 3.340 3.590 ;
        RECT  3.180 3.390 3.340 4.480 ;
        RECT  3.180 4.320 4.520 4.480 ;
        RECT  2.510 0.320 4.780 0.480 ;
        RECT  2.510 0.320 2.710 1.220 ;
        RECT  2.510 1.060 3.420 1.220 ;
        RECT  3.220 1.060 3.420 1.740 ;
        RECT  3.860 2.760 4.060 3.120 ;
        RECT  5.220 2.880 5.500 3.120 ;
        RECT  3.860 2.960 5.500 3.120 ;
        RECT  3.180 2.880 3.660 3.040 ;
        RECT  3.500 2.880 3.660 3.850 ;
        RECT  3.500 3.650 5.600 3.850 ;
        RECT  3.820 3.650 4.100 4.160 ;
        RECT  5.740 2.990 5.940 3.440 ;
        RECT  4.160 3.280 5.940 3.440 ;
        RECT  5.780 2.990 5.940 4.420 ;
        RECT  5.780 4.220 6.180 4.420 ;
        RECT  3.100 0.640 3.740 0.800 ;
        RECT  3.580 0.640 3.740 1.280 ;
        RECT  3.580 1.120 6.240 1.280 ;
        RECT  3.740 1.120 3.940 1.740 ;
        RECT  3.940 0.640 4.220 0.960 ;
        RECT  7.390 0.680 7.670 0.960 ;
        RECT  3.940 0.800 7.670 0.960 ;
        RECT  4.340 1.440 7.700 1.600 ;
        RECT  7.420 1.440 7.700 1.720 ;
        RECT  4.340 1.440 4.540 1.750 ;
        RECT  5.380 1.760 7.120 1.920 ;
        RECT  6.960 1.760 7.120 2.100 ;
        RECT  6.960 1.940 7.900 2.100 ;
        RECT  7.060 0.300 7.910 0.500 ;
        RECT  5.700 0.480 7.220 0.640 ;
        LAYER VTPH ;
        RECT  1.790 1.140 2.630 3.640 ;
        RECT  0.000 1.140 0.850 3.660 ;
        RECT  1.790 1.160 7.150 3.640 ;
        RECT  4.470 1.140 7.150 3.640 ;
        RECT  0.000 1.190 1.900 3.660 ;
        RECT  4.880 1.200 8.400 3.660 ;
        LAYER VTNH ;
        RECT  1.900 3.640 4.880 4.800 ;
        RECT  0.000 3.660 8.400 4.800 ;
        RECT  0.000 0.000 8.400 1.140 ;
        RECT  2.630 0.000 4.470 1.160 ;
        RECT  0.850 0.000 1.790 1.190 ;
        RECT  7.150 0.000 8.400 1.200 ;
    END
END SDFQRM4HM

MACRO SDFQRM2HM
    CLASS CORE ;
    FOREIGN SDFQRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        ANTENNAGATEAREA 0.102  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.518  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.860 0.930 2.060 1.130 ;
        LAYER ME2 ;
        RECT  1.700 0.830 2.060 1.230 ;
        LAYER ME1 ;
        RECT  1.780 0.900 2.150 1.220 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        ANTENNAGATEAREA 0.062  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.833  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.800 1.060 3.000 1.260 ;
        LAYER ME2 ;
        RECT  2.800 0.840 3.100 1.360 ;
        LAYER ME1 ;
        RECT  2.800 0.900 3.040 1.360 ;
        END
    END CK
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        ANTENNAGATEAREA 0.115  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.250  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.100 1.080 10.300 1.280 ;
        LAYER ME2 ;
        RECT  10.100 0.840 10.300 1.380 ;
        LAYER ME1 ;
        RECT  9.910 1.080 10.430 1.280 ;
        END
    END RB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.660 0.420 11.900 2.100 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.140 1.290 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.290 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  11.040 2.080 11.320 2.540 ;
        RECT  10.020 1.840 10.220 2.540 ;
        RECT  7.240 1.860 7.520 2.540 ;
        RECT  6.300 1.440 6.500 2.540 ;
        RECT  2.660 2.020 2.860 2.540 ;
        RECT  0.660 1.840 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  11.080 -0.140 11.360 0.540 ;
        RECT  9.700 -0.140 9.980 0.540 ;
        RECT  7.520 -0.140 7.680 0.690 ;
        RECT  2.600 -0.140 2.760 0.420 ;
        RECT  0.620 -0.140 0.900 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.460 0.380 0.660 ;
        RECT  0.100 0.460 0.260 1.920 ;
        RECT  1.400 1.380 2.560 1.540 ;
        RECT  2.360 0.900 2.560 1.540 ;
        RECT  1.400 1.180 1.600 1.680 ;
        RECT  0.100 1.520 1.600 1.680 ;
        RECT  0.100 1.520 0.340 1.920 ;
        RECT  3.240 0.620 3.520 0.840 ;
        RECT  3.340 0.620 3.520 1.300 ;
        RECT  3.340 1.100 4.100 1.300 ;
        RECT  3.340 0.620 3.500 1.780 ;
        RECT  4.160 0.620 4.440 0.840 ;
        RECT  4.260 0.620 4.440 1.190 ;
        RECT  4.260 1.030 4.820 1.190 ;
        RECT  4.260 0.620 4.420 1.760 ;
        RECT  2.920 0.300 4.860 0.460 ;
        RECT  1.540 0.400 2.280 0.560 ;
        RECT  2.100 0.400 2.280 0.740 ;
        RECT  4.700 0.300 4.860 0.700 ;
        RECT  2.920 0.300 3.080 0.740 ;
        RECT  2.100 0.580 3.080 0.740 ;
        RECT  2.140 1.700 3.180 1.860 ;
        RECT  3.020 1.700 3.180 2.100 ;
        RECT  1.540 1.860 2.300 2.020 ;
        RECT  4.720 1.520 4.920 2.100 ;
        RECT  3.020 1.940 4.920 2.100 ;
        RECT  5.220 0.440 5.380 1.720 ;
        RECT  5.220 0.660 7.040 0.820 ;
        RECT  6.840 0.660 7.040 0.940 ;
        RECT  5.220 0.660 5.420 1.720 ;
        RECT  5.880 1.100 6.820 1.260 ;
        RECT  5.880 1.100 6.080 1.380 ;
        RECT  6.660 1.100 6.820 1.680 ;
        RECT  8.160 0.620 8.360 1.680 ;
        RECT  6.660 1.520 8.360 1.680 ;
        RECT  7.880 1.520 8.080 2.080 ;
        RECT  7.840 0.300 9.360 0.460 ;
        RECT  5.540 0.300 7.360 0.500 ;
        RECT  7.200 0.300 7.360 1.010 ;
        RECT  7.840 0.300 8.000 1.010 ;
        RECT  7.200 0.850 8.000 1.010 ;
        RECT  8.520 0.300 8.680 1.340 ;
        RECT  9.200 0.300 9.360 1.580 ;
        RECT  9.200 1.380 9.540 1.580 ;
        RECT  9.700 1.440 10.980 1.600 ;
        RECT  8.840 0.630 9.040 1.920 ;
        RECT  8.840 1.760 9.860 1.920 ;
        RECT  9.700 1.440 9.860 1.920 ;
        RECT  8.360 1.840 9.030 2.040 ;
        RECT  10.620 0.300 10.780 0.860 ;
        RECT  9.540 0.700 11.480 0.860 ;
        RECT  9.540 0.700 9.700 1.180 ;
        RECT  11.320 0.700 11.480 1.920 ;
        RECT  10.520 1.760 11.480 1.920 ;
        RECT  10.520 1.760 10.720 2.100 ;
        LAYER VTPH ;
        RECT  1.590 1.120 2.450 2.400 ;
        RECT  0.000 1.140 7.250 2.400 ;
        RECT  9.620 1.140 12.000 2.400 ;
        RECT  0.000 1.210 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.120 ;
        RECT  0.000 0.000 1.590 1.140 ;
        RECT  2.450 0.000 12.000 1.140 ;
        RECT  7.250 0.000 9.620 1.210 ;
    END
END SDFQRM2HM

MACRO SDFQRM1HM
    CLASS CORE ;
    FOREIGN SDFQRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        ANTENNAGATEAREA 0.102  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.518  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.860 0.930 2.060 1.130 ;
        LAYER ME2 ;
        RECT  1.700 0.830 2.060 1.230 ;
        LAYER ME1 ;
        RECT  1.780 0.900 2.150 1.220 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        ANTENNAGATEAREA 0.062  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.833  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.800 1.060 3.000 1.260 ;
        LAYER ME2 ;
        RECT  2.800 0.840 3.100 1.360 ;
        LAYER ME1 ;
        RECT  2.800 0.900 3.040 1.360 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.660 0.380 11.900 2.000 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.140 1.290 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.290 ;
        END
    END SE
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        ANTENNAGATEAREA 0.115  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.250  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.100 1.080 10.300 1.280 ;
        LAYER ME2 ;
        RECT  10.100 0.840 10.300 1.380 ;
        LAYER ME1 ;
        RECT  9.910 1.080 10.430 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  11.040 2.080 11.320 2.540 ;
        RECT  10.020 1.840 10.220 2.540 ;
        RECT  7.240 1.860 7.520 2.540 ;
        RECT  6.300 1.440 6.500 2.540 ;
        RECT  2.660 2.020 2.860 2.540 ;
        RECT  0.660 1.840 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  11.080 -0.140 11.360 0.540 ;
        RECT  9.700 -0.140 9.980 0.540 ;
        RECT  7.520 -0.140 7.680 0.690 ;
        RECT  2.600 -0.140 2.760 0.420 ;
        RECT  0.620 -0.140 0.900 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.460 0.380 0.660 ;
        RECT  0.100 0.460 0.260 1.920 ;
        RECT  1.400 1.380 2.560 1.540 ;
        RECT  2.360 0.900 2.560 1.540 ;
        RECT  1.400 1.180 1.600 1.680 ;
        RECT  0.100 1.520 1.600 1.680 ;
        RECT  0.100 1.520 0.340 1.920 ;
        RECT  3.240 0.620 3.520 0.840 ;
        RECT  3.340 0.620 3.520 1.300 ;
        RECT  3.340 1.100 4.100 1.300 ;
        RECT  3.340 0.620 3.500 1.780 ;
        RECT  4.160 0.620 4.440 0.840 ;
        RECT  4.260 0.620 4.440 1.190 ;
        RECT  4.260 1.030 4.820 1.190 ;
        RECT  4.260 0.620 4.420 1.760 ;
        RECT  2.920 0.300 4.860 0.460 ;
        RECT  1.540 0.400 2.280 0.560 ;
        RECT  2.100 0.400 2.280 0.740 ;
        RECT  4.700 0.300 4.860 0.700 ;
        RECT  2.920 0.300 3.080 0.740 ;
        RECT  2.100 0.580 3.080 0.740 ;
        RECT  2.140 1.700 3.180 1.860 ;
        RECT  3.020 1.700 3.180 2.100 ;
        RECT  1.540 1.860 2.300 2.020 ;
        RECT  4.720 1.520 4.920 2.100 ;
        RECT  3.020 1.940 4.920 2.100 ;
        RECT  5.220 0.440 5.380 1.720 ;
        RECT  5.220 0.660 7.040 0.820 ;
        RECT  6.840 0.660 7.040 0.940 ;
        RECT  5.220 0.660 5.420 1.720 ;
        RECT  5.880 1.100 6.820 1.260 ;
        RECT  5.880 1.100 6.080 1.380 ;
        RECT  6.660 1.100 6.820 1.680 ;
        RECT  8.160 0.620 8.360 1.680 ;
        RECT  6.660 1.520 8.360 1.680 ;
        RECT  7.880 1.520 8.080 2.080 ;
        RECT  7.840 0.300 9.360 0.460 ;
        RECT  5.540 0.300 7.360 0.500 ;
        RECT  7.200 0.300 7.360 1.010 ;
        RECT  7.840 0.300 8.000 1.010 ;
        RECT  7.200 0.850 8.000 1.010 ;
        RECT  8.520 0.300 8.680 1.340 ;
        RECT  9.200 0.300 9.360 1.580 ;
        RECT  9.200 1.380 9.540 1.580 ;
        RECT  9.700 1.440 10.980 1.600 ;
        RECT  8.840 0.630 9.040 1.920 ;
        RECT  8.840 1.760 9.860 1.920 ;
        RECT  9.700 1.440 9.860 1.920 ;
        RECT  8.360 1.840 9.030 2.040 ;
        RECT  10.620 0.300 10.780 0.860 ;
        RECT  9.540 0.700 11.480 0.860 ;
        RECT  9.540 0.700 9.700 1.180 ;
        RECT  11.320 0.700 11.480 1.920 ;
        RECT  10.520 1.760 11.480 1.920 ;
        RECT  10.520 1.760 10.720 2.100 ;
        LAYER VTPH ;
        RECT  1.590 1.120 2.450 2.400 ;
        RECT  0.000 1.140 7.250 2.400 ;
        RECT  9.620 1.140 12.000 2.400 ;
        RECT  0.000 1.210 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.120 ;
        RECT  0.000 0.000 1.590 1.140 ;
        RECT  2.450 0.000 12.000 1.140 ;
        RECT  7.250 0.000 9.620 1.210 ;
    END
END SDFQRM1HM

MACRO SDFQM8HM
    CLASS CORE ;
    FOREIGN SDFQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.564  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.610 1.090 2.810 1.290 ;
        LAYER ME2 ;
        RECT  2.500 0.900 2.810 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.040 2.910 1.340 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.853  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.160 1.170 3.360 1.370 ;
        LAYER ME2 ;
        RECT  3.130 0.900 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.070 1.060 3.440 1.480 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.900 0.730 12.170 2.100 ;
        RECT  11.910 0.380 12.170 2.100 ;
        RECT  10.890 1.370 12.170 1.560 ;
        RECT  11.700 0.730 12.170 1.560 ;
        RECT  10.890 0.730 12.170 0.890 ;
        RECT  10.890 1.370 11.120 2.100 ;
        RECT  10.890 0.420 11.110 0.890 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.450 0.710 1.640 0.880 ;
        RECT  0.450 0.710 0.700 1.190 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.839  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.900 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.050 1.200 1.380 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  12.460 1.460 12.660 2.540 ;
        RECT  11.420 1.840 11.620 2.540 ;
        RECT  9.480 2.020 9.680 2.540 ;
        RECT  7.150 1.860 7.430 2.540 ;
        RECT  4.320 1.970 4.480 2.540 ;
        RECT  2.950 1.980 3.110 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  12.460 -0.140 12.660 0.710 ;
        RECT  11.380 -0.140 11.660 0.520 ;
        RECT  9.270 -0.140 9.560 0.400 ;
        RECT  7.150 -0.140 7.370 0.400 ;
        RECT  4.400 -0.140 4.560 0.420 ;
        RECT  2.940 -0.140 3.140 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.560 ;
        RECT  0.100 0.300 0.260 2.100 ;
        RECT  1.820 0.820 2.020 1.700 ;
        RECT  0.100 1.540 2.020 1.700 ;
        RECT  0.100 1.540 0.340 2.100 ;
        RECT  2.180 0.620 2.460 0.840 ;
        RECT  2.180 0.620 2.340 1.700 ;
        RECT  2.180 1.500 2.460 1.700 ;
        RECT  3.620 0.620 3.900 1.200 ;
        RECT  3.620 1.000 4.690 1.200 ;
        RECT  3.620 0.620 3.840 1.760 ;
        RECT  5.040 0.620 5.320 1.720 ;
        RECT  5.040 1.260 5.500 1.720 ;
        RECT  4.960 1.440 5.500 1.720 ;
        RECT  4.000 1.550 4.800 1.710 ;
        RECT  2.620 1.660 3.440 1.820 ;
        RECT  3.280 1.660 3.440 2.100 ;
        RECT  4.640 1.550 4.800 2.100 ;
        RECT  2.620 1.660 2.780 2.020 ;
        RECT  1.500 1.860 2.780 2.020 ;
        RECT  4.000 1.550 4.160 2.100 ;
        RECT  3.280 1.940 4.160 2.100 ;
        RECT  5.300 1.900 5.580 2.100 ;
        RECT  4.640 1.940 5.580 2.100 ;
        RECT  1.460 0.300 2.780 0.460 ;
        RECT  3.300 0.300 4.220 0.460 ;
        RECT  4.720 0.300 5.840 0.460 ;
        RECT  1.460 0.300 1.830 0.500 ;
        RECT  5.520 0.300 5.840 0.560 ;
        RECT  4.060 0.300 4.220 0.740 ;
        RECT  2.620 0.300 2.780 0.880 ;
        RECT  4.720 0.300 4.880 0.740 ;
        RECT  4.060 0.580 4.880 0.740 ;
        RECT  3.300 0.300 3.460 0.880 ;
        RECT  2.620 0.720 3.460 0.880 ;
        RECT  5.480 0.760 5.900 1.040 ;
        RECT  5.740 0.760 5.900 2.100 ;
        RECT  5.740 1.940 6.720 2.100 ;
        RECT  6.060 0.920 7.580 1.120 ;
        RECT  6.060 0.300 6.260 1.780 ;
        RECT  6.770 1.300 8.080 1.520 ;
        RECT  7.860 0.620 8.080 1.850 ;
        RECT  7.770 1.300 8.080 1.850 ;
        RECT  7.530 0.300 8.890 0.460 ;
        RECT  7.530 0.300 7.690 0.760 ;
        RECT  6.450 0.560 7.690 0.760 ;
        RECT  8.730 0.300 8.890 1.780 ;
        RECT  8.720 1.560 9.000 1.780 ;
        RECT  8.290 0.620 8.540 0.900 ;
        RECT  9.520 0.980 9.740 1.860 ;
        RECT  9.160 1.700 9.740 1.860 ;
        RECT  8.290 0.620 8.450 2.100 ;
        RECT  9.160 1.700 9.320 2.100 ;
        RECT  8.290 1.940 9.320 2.100 ;
        RECT  9.100 0.620 10.180 0.820 ;
        RECT  9.920 0.620 10.180 1.210 ;
        RECT  9.920 1.050 11.530 1.210 ;
        RECT  9.100 0.620 9.300 1.360 ;
        RECT  9.920 0.620 10.120 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.470 2.400 ;
        RECT  8.910 1.140 12.800 2.400 ;
        RECT  0.000 1.200 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
        RECT  7.470 0.000 8.910 1.200 ;
    END
END SDFQM8HM

MACRO SDFQM4HM
    CLASS CORE ;
    FOREIGN SDFQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.349  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.160 1.170 3.360 1.370 ;
        LAYER ME2 ;
        RECT  3.130 0.900 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.070 1.060 3.440 1.480 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.564  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.610 1.090 2.810 1.290 ;
        LAYER ME2 ;
        RECT  2.500 0.900 2.810 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.040 2.910 1.340 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.000 1.370 11.900 1.560 ;
        RECT  11.700 0.730 11.900 1.560 ;
        RECT  11.000 0.730 11.900 0.890 ;
        RECT  11.000 1.370 11.320 2.100 ;
        RECT  11.000 0.370 11.320 0.890 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.450 0.710 1.640 0.880 ;
        RECT  0.450 0.710 0.700 1.190 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.839  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.900 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.050 1.200 1.380 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  11.580 1.840 11.780 2.540 ;
        RECT  10.560 1.510 10.760 2.540 ;
        RECT  9.480 1.710 9.680 2.540 ;
        RECT  7.150 1.860 7.430 2.540 ;
        RECT  4.320 1.970 4.480 2.540 ;
        RECT  2.950 1.980 3.110 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  11.540 -0.140 11.820 0.520 ;
        RECT  10.540 -0.140 10.740 0.840 ;
        RECT  9.270 -0.140 9.560 0.400 ;
        RECT  7.150 -0.140 7.370 0.400 ;
        RECT  4.400 -0.140 4.560 0.420 ;
        RECT  2.940 -0.140 3.140 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.560 ;
        RECT  0.100 0.300 0.260 2.100 ;
        RECT  1.820 0.820 2.020 1.700 ;
        RECT  0.100 1.540 2.020 1.700 ;
        RECT  0.100 1.540 0.340 2.100 ;
        RECT  2.180 0.620 2.460 0.840 ;
        RECT  2.180 0.620 2.340 1.700 ;
        RECT  2.180 1.500 2.460 1.700 ;
        RECT  3.620 0.620 3.900 1.200 ;
        RECT  3.620 1.000 4.690 1.200 ;
        RECT  3.620 0.620 3.840 1.760 ;
        RECT  5.040 0.620 5.320 1.720 ;
        RECT  5.040 1.260 5.500 1.720 ;
        RECT  4.960 1.440 5.500 1.720 ;
        RECT  4.000 1.550 4.800 1.710 ;
        RECT  2.620 1.660 3.440 1.820 ;
        RECT  4.640 1.550 4.800 2.100 ;
        RECT  3.280 1.660 3.440 2.100 ;
        RECT  2.620 1.660 2.780 2.020 ;
        RECT  1.500 1.860 2.780 2.020 ;
        RECT  4.000 1.550 4.160 2.100 ;
        RECT  3.280 1.940 4.160 2.100 ;
        RECT  4.640 1.900 5.580 2.100 ;
        RECT  1.460 0.300 2.780 0.460 ;
        RECT  3.300 0.300 4.220 0.460 ;
        RECT  4.720 0.300 5.840 0.460 ;
        RECT  1.460 0.300 1.830 0.500 ;
        RECT  5.520 0.300 5.840 0.560 ;
        RECT  4.060 0.300 4.220 0.740 ;
        RECT  2.620 0.300 2.780 0.880 ;
        RECT  4.720 0.300 4.880 0.740 ;
        RECT  4.060 0.580 4.880 0.740 ;
        RECT  3.300 0.300 3.460 0.880 ;
        RECT  2.620 0.720 3.460 0.880 ;
        RECT  5.480 0.760 5.900 1.040 ;
        RECT  5.740 0.760 5.900 2.100 ;
        RECT  5.740 1.940 6.720 2.100 ;
        RECT  6.060 0.920 7.580 1.120 ;
        RECT  6.060 0.300 6.260 1.780 ;
        RECT  6.770 1.300 8.080 1.520 ;
        RECT  7.860 0.620 8.080 1.850 ;
        RECT  7.770 1.300 8.080 1.850 ;
        RECT  7.530 0.300 8.890 0.460 ;
        RECT  7.530 0.300 7.690 0.760 ;
        RECT  6.450 0.560 7.690 0.760 ;
        RECT  8.720 0.300 8.890 1.780 ;
        RECT  8.720 1.560 9.000 1.780 ;
        RECT  9.520 0.980 9.740 1.540 ;
        RECT  9.160 1.380 9.740 1.540 ;
        RECT  8.290 0.620 8.540 2.100 ;
        RECT  9.160 1.380 9.320 2.100 ;
        RECT  8.290 1.940 9.320 2.100 ;
        RECT  9.100 0.620 10.300 0.820 ;
        RECT  10.040 0.620 10.300 1.210 ;
        RECT  10.040 1.050 11.180 1.210 ;
        RECT  9.100 0.620 9.300 1.220 ;
        RECT  10.040 0.620 10.240 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.470 2.400 ;
        RECT  8.910 1.140 12.000 2.400 ;
        RECT  0.000 1.200 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.140 ;
        RECT  7.470 0.000 8.910 1.200 ;
    END
END SDFQM4HM

MACRO SDFQM2HM
    CLASS CORE ;
    FOREIGN SDFQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.564  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.610 1.090 2.810 1.290 ;
        LAYER ME2 ;
        RECT  2.500 0.900 2.810 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.040 2.910 1.340 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.349  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.160 1.170 3.360 1.370 ;
        LAYER ME2 ;
        RECT  3.130 0.900 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.070 1.060 3.440 1.480 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.800 0.370 11.100 2.100 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.450 0.710 1.640 0.880 ;
        RECT  0.450 0.710 0.700 1.190 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.839  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.900 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.050 1.200 1.380 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.260 2.080 10.540 2.540 ;
        RECT  9.450 1.710 9.650 2.540 ;
        RECT  7.150 1.860 7.430 2.540 ;
        RECT  4.320 1.970 4.480 2.540 ;
        RECT  2.950 1.980 3.110 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.340 -0.140 10.540 0.560 ;
        RECT  9.140 -0.140 9.430 0.400 ;
        RECT  7.150 -0.140 7.370 0.400 ;
        RECT  4.400 -0.140 4.560 0.420 ;
        RECT  2.940 -0.140 3.140 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.560 ;
        RECT  0.100 0.300 0.260 2.100 ;
        RECT  1.820 0.820 2.020 1.700 ;
        RECT  0.100 1.540 2.020 1.700 ;
        RECT  0.100 1.540 0.340 2.100 ;
        RECT  2.180 0.620 2.460 0.840 ;
        RECT  2.180 0.620 2.340 1.700 ;
        RECT  2.180 1.500 2.460 1.700 ;
        RECT  3.620 0.620 3.900 1.200 ;
        RECT  3.620 1.000 4.690 1.200 ;
        RECT  3.620 0.620 3.840 1.760 ;
        RECT  5.040 0.620 5.320 1.720 ;
        RECT  5.040 1.260 5.500 1.720 ;
        RECT  4.960 1.440 5.500 1.720 ;
        RECT  4.000 1.550 4.800 1.710 ;
        RECT  2.620 1.660 3.440 1.820 ;
        RECT  4.640 1.550 4.800 2.100 ;
        RECT  3.280 1.660 3.440 2.100 ;
        RECT  2.620 1.660 2.780 2.020 ;
        RECT  1.500 1.860 2.780 2.020 ;
        RECT  4.000 1.550 4.160 2.100 ;
        RECT  3.280 1.940 4.160 2.100 ;
        RECT  4.640 1.900 5.580 2.100 ;
        RECT  1.460 0.300 2.780 0.460 ;
        RECT  3.300 0.300 4.220 0.460 ;
        RECT  4.720 0.300 5.840 0.460 ;
        RECT  1.460 0.300 1.830 0.500 ;
        RECT  5.520 0.300 5.840 0.560 ;
        RECT  4.060 0.300 4.220 0.740 ;
        RECT  2.620 0.300 2.780 0.880 ;
        RECT  4.720 0.300 4.880 0.740 ;
        RECT  4.060 0.580 4.880 0.740 ;
        RECT  3.300 0.300 3.460 0.880 ;
        RECT  2.620 0.720 3.460 0.880 ;
        RECT  5.480 0.760 5.900 1.040 ;
        RECT  5.740 0.760 5.900 2.100 ;
        RECT  5.740 1.940 6.720 2.100 ;
        RECT  6.060 0.920 7.580 1.120 ;
        RECT  6.060 0.300 6.260 1.780 ;
        RECT  6.770 1.300 8.080 1.520 ;
        RECT  7.860 0.620 8.080 1.850 ;
        RECT  7.770 1.300 8.080 1.850 ;
        RECT  7.530 0.300 8.930 0.460 ;
        RECT  7.530 0.300 7.690 0.760 ;
        RECT  6.450 0.560 7.690 0.760 ;
        RECT  8.770 0.300 8.930 1.780 ;
        RECT  8.690 1.560 8.970 1.780 ;
        RECT  8.290 0.620 8.540 0.900 ;
        RECT  9.510 0.980 9.750 1.540 ;
        RECT  9.130 1.380 9.750 1.540 ;
        RECT  8.290 0.620 8.450 2.100 ;
        RECT  9.130 1.380 9.290 2.100 ;
        RECT  8.290 1.940 9.290 2.100 ;
        RECT  9.090 0.620 10.190 0.820 ;
        RECT  9.990 0.620 10.190 1.270 ;
        RECT  9.090 0.620 9.290 1.220 ;
        RECT  9.990 0.990 10.630 1.270 ;
        RECT  9.990 0.620 10.150 1.760 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.470 2.400 ;
        RECT  8.900 1.140 11.200 2.400 ;
        RECT  0.000 1.200 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
        RECT  7.470 0.000 8.900 1.200 ;
    END
END SDFQM2HM

MACRO SDFQM1HM
    CLASS CORE ;
    FOREIGN SDFQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER ME1  ;
        ANTENNAGATEAREA 0.160  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.737  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.300 1.110 0.500 1.310 ;
        LAYER ME2 ;
        RECT  0.300 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.040 0.600 1.380 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        ANTENNAGATEAREA 0.038  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.833  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.110 1.100 1.310 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.800 1.040 1.260 1.380 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.760 3.200 1.230 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.980 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.080 0.460 10.300 1.830 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.420 2.080 9.740 2.540 ;
        RECT  6.500 2.080 6.780 2.540 ;
        RECT  2.800 2.020 3.020 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.480 -0.140 9.680 0.710 ;
        RECT  6.340 -0.140 6.540 0.380 ;
        RECT  4.400 -0.140 4.680 0.320 ;
        RECT  2.660 -0.140 2.940 0.500 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.300 2.380 0.460 ;
        RECT  2.220 0.300 2.380 0.820 ;
        RECT  0.160 0.470 0.320 0.880 ;
        RECT  2.220 0.660 2.700 0.820 ;
        RECT  0.160 0.720 1.580 0.880 ;
        RECT  2.480 0.660 2.700 1.050 ;
        RECT  1.420 0.300 1.580 1.700 ;
        RECT  0.160 1.540 1.580 1.700 ;
        RECT  0.160 1.540 0.320 1.990 ;
        RECT  3.360 0.350 3.680 0.630 ;
        RECT  3.520 0.350 3.680 1.710 ;
        RECT  1.740 0.620 2.020 0.820 ;
        RECT  4.600 1.120 4.900 1.320 ;
        RECT  2.460 1.560 3.350 1.720 ;
        RECT  1.740 0.620 1.900 2.040 ;
        RECT  3.190 1.560 3.350 2.100 ;
        RECT  2.460 1.560 2.620 2.040 ;
        RECT  1.740 1.880 2.620 2.040 ;
        RECT  4.600 1.120 4.760 2.100 ;
        RECT  3.190 1.940 4.760 2.100 ;
        RECT  5.480 0.620 5.760 1.280 ;
        RECT  5.480 1.000 6.960 1.280 ;
        RECT  5.480 0.620 5.700 1.780 ;
        RECT  5.380 1.440 5.700 1.780 ;
        RECT  7.090 0.620 7.420 0.900 ;
        RECT  7.260 0.620 7.420 1.780 ;
        RECT  6.240 1.440 7.460 1.600 ;
        RECT  7.260 1.440 7.460 1.780 ;
        RECT  4.200 0.800 5.320 0.960 ;
        RECT  5.150 0.700 5.320 1.060 ;
        RECT  4.200 0.800 4.420 1.080 ;
        RECT  5.860 1.760 7.100 1.920 ;
        RECT  5.060 0.800 5.220 2.100 ;
        RECT  6.940 1.760 7.100 2.100 ;
        RECT  5.860 1.500 6.080 2.100 ;
        RECT  5.060 1.940 6.080 2.100 ;
        RECT  6.940 1.940 7.680 2.100 ;
        RECT  4.840 0.300 6.180 0.460 ;
        RECT  6.700 0.300 8.320 0.460 ;
        RECT  3.880 0.300 4.080 0.640 ;
        RECT  5.920 0.300 6.180 0.700 ;
        RECT  4.840 0.300 5.000 0.640 ;
        RECT  3.880 0.480 5.000 0.640 ;
        RECT  6.700 0.300 6.860 0.700 ;
        RECT  5.920 0.540 6.860 0.700 ;
        RECT  8.160 0.300 8.320 1.720 ;
        RECT  3.880 0.300 4.040 1.700 ;
        RECT  3.880 1.500 4.220 1.700 ;
        RECT  8.160 1.360 8.380 1.720 ;
        RECT  8.780 0.530 9.150 0.730 ;
        RECT  8.780 0.530 8.940 1.600 ;
        RECT  8.780 1.400 9.140 1.600 ;
        RECT  7.610 0.620 8.000 0.900 ;
        RECT  9.300 0.990 9.810 1.200 ;
        RECT  9.300 0.990 9.460 1.920 ;
        RECT  8.540 1.760 9.460 1.920 ;
        RECT  7.840 0.620 8.000 2.100 ;
        RECT  8.540 1.760 8.700 2.100 ;
        RECT  7.840 1.940 8.700 2.100 ;
        LAYER VTPH ;
        RECT  2.190 1.090 4.740 2.400 ;
        RECT  8.680 1.050 9.850 2.400 ;
        RECT  0.000 1.140 5.630 2.400 ;
        RECT  8.030 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.050 ;
        RECT  0.000 0.000 8.680 1.090 ;
        RECT  0.000 0.000 2.190 1.140 ;
        RECT  4.740 0.000 8.680 1.140 ;
        RECT  9.850 0.000 10.400 1.140 ;
        RECT  5.630 0.000 8.030 1.200 ;
    END
END SDFQM1HM

MACRO SDFMQM8HM
    CLASS CORE ;
    FOREIGN SDFMQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.706  LAYER ME1  ;
        ANTENNADIFFAREA 1.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.770 0.400 9.100 1.720 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  6.010 2.260 6.290 2.720 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.300 -0.140 9.560 0.750 ;
        RECT  8.280 -0.140 8.480 0.700 ;
        RECT  7.240 -0.140 7.460 0.610 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 10.000 4.940 ;
        RECT  9.300 3.970 9.540 4.940 ;
        RECT  8.300 4.240 8.500 4.940 ;
        RECT  6.020 4.480 6.300 4.940 ;
        RECT  3.630 4.320 3.830 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.880 0.320 3.240 ;
        RECT  0.100 2.880 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.130 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.290 ;
        RECT  6.750 3.770 7.100 4.000 ;
        RECT  4.750 3.840 7.100 4.000 ;
        RECT  3.050 4.000 4.230 4.160 ;
        RECT  3.050 4.000 3.390 4.290 ;
        RECT  4.070 4.000 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.810 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.600 2.700 7.810 4.150 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.420 3.360 ;
        RECT  4.850 3.200 7.420 3.360 ;
        RECT  8.430 3.580 8.650 4.080 ;
        RECT  7.970 3.920 8.650 4.080 ;
        RECT  5.070 4.160 7.420 4.320 ;
        RECT  7.260 3.060 7.420 4.500 ;
        RECT  7.010 4.160 7.420 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.970 3.920 8.130 4.500 ;
        RECT  7.010 4.340 8.130 4.500 ;
        RECT  8.750 3.140 9.050 3.360 ;
        RECT  8.810 3.140 9.050 4.470 ;
        RECT  8.010 2.820 9.420 2.980 ;
        RECT  9.240 2.820 9.420 3.810 ;
        RECT  8.010 2.820 8.210 3.630 ;
        RECT  9.240 3.560 9.730 3.810 ;
        RECT  9.310 0.990 9.830 1.240 ;
        RECT  7.780 0.560 7.980 2.060 ;
        RECT  7.660 1.690 7.980 2.060 ;
        RECT  9.310 0.990 9.470 2.060 ;
        RECT  7.660 1.900 9.470 2.060 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 10.000 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 10.000 3.660 ;
        RECT  4.820 1.180 10.000 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 10.000 4.800 ;
        RECT  0.000 0.000 10.000 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 10.000 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMQM8HM

MACRO SDFMQM4HM
    CLASS CORE ;
    FOREIGN SDFMQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.738  LAYER ME1  ;
        ANTENNADIFFAREA 0.896  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.780 0.550 9.160 1.570 ;
        RECT  8.780 0.550 9.060 1.720 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  6.010 2.260 6.290 2.720 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.290 -0.140 8.490 0.710 ;
        RECT  7.270 -0.140 7.490 0.440 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  8.310 4.240 8.510 4.940 ;
        RECT  6.020 4.480 6.300 4.940 ;
        RECT  3.610 4.480 3.890 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.950 0.320 3.300 ;
        RECT  0.100 2.950 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.240 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.250 ;
        RECT  6.750 3.770 7.100 4.000 ;
        RECT  4.750 3.840 7.100 4.000 ;
        RECT  3.050 3.970 4.230 4.250 ;
        RECT  4.070 3.970 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.810 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.600 2.700 7.810 4.150 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.420 3.360 ;
        RECT  4.850 3.200 7.420 3.360 ;
        RECT  8.430 3.580 8.660 4.080 ;
        RECT  7.970 3.920 8.660 4.080 ;
        RECT  5.070 4.160 7.420 4.320 ;
        RECT  7.260 3.060 7.420 4.500 ;
        RECT  7.010 4.160 7.420 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.970 3.920 8.130 4.500 ;
        RECT  7.010 4.340 8.130 4.500 ;
        RECT  8.760 3.140 9.060 3.360 ;
        RECT  8.820 3.140 9.060 4.260 ;
        RECT  8.010 2.820 9.490 2.980 ;
        RECT  9.270 2.820 9.490 3.100 ;
        RECT  8.010 2.820 8.210 3.630 ;
        RECT  7.780 0.560 7.980 2.060 ;
        RECT  7.660 1.480 7.980 2.060 ;
        RECT  9.210 1.780 9.490 2.060 ;
        RECT  7.660 1.900 9.490 2.060 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 9.600 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 9.600 3.660 ;
        RECT  4.820 1.180 9.600 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 9.600 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMQM4HM

MACRO SDFMQM2HM
    CLASS CORE ;
    FOREIGN SDFMQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.371  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.760 3.080 9.100 3.960 ;
        RECT  8.570 4.130 8.920 4.370 ;
        RECT  8.760 3.080 8.920 4.370 ;
        RECT  8.640 3.080 9.100 3.360 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.440 -0.140 8.650 0.870 ;
        RECT  7.270 -0.140 7.490 0.440 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 9.200 4.940 ;
        RECT  8.150 4.240 8.350 4.940 ;
        RECT  5.900 4.480 6.180 4.940 ;
        RECT  3.610 4.480 3.890 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.950 0.320 3.300 ;
        RECT  0.100 2.950 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.240 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.250 ;
        RECT  4.750 3.840 6.930 4.000 ;
        RECT  3.050 3.970 4.230 4.250 ;
        RECT  4.070 3.970 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.610 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.410 2.700 7.610 4.160 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.250 3.360 ;
        RECT  4.850 3.200 7.250 3.360 ;
        RECT  8.360 3.580 8.580 3.950 ;
        RECT  7.830 3.790 8.580 3.950 ;
        RECT  5.070 4.160 7.250 4.320 ;
        RECT  7.090 3.060 7.250 4.500 ;
        RECT  6.780 4.160 7.250 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.830 3.790 7.990 4.500 ;
        RECT  6.780 4.340 7.990 4.500 ;
        RECT  7.850 0.560 8.050 2.050 ;
        RECT  7.690 1.770 8.960 2.050 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 9.200 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 9.200 3.660 ;
        RECT  4.820 1.180 9.200 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 9.200 4.800 ;
        RECT  0.000 0.000 9.200 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 9.200 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMQM2HM

MACRO SDFMQM1HM
    CLASS CORE ;
    FOREIGN SDFMQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.760 3.390 9.100 3.960 ;
        RECT  8.570 4.260 8.920 4.500 ;
        RECT  8.760 3.080 8.920 4.500 ;
        RECT  8.640 3.080 8.920 3.360 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.440 -0.140 8.650 0.870 ;
        RECT  7.270 -0.140 7.490 0.440 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 9.200 4.940 ;
        RECT  8.150 4.240 8.350 4.940 ;
        RECT  5.900 4.480 6.180 4.940 ;
        RECT  3.610 4.480 3.890 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.950 0.320 3.300 ;
        RECT  0.100 2.950 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.240 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.250 ;
        RECT  4.750 3.840 6.930 4.000 ;
        RECT  3.050 3.970 4.230 4.250 ;
        RECT  4.070 3.970 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.610 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.410 2.700 7.610 4.160 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.250 3.360 ;
        RECT  4.850 3.200 7.250 3.360 ;
        RECT  8.360 3.580 8.580 3.950 ;
        RECT  7.830 3.790 8.580 3.950 ;
        RECT  5.070 4.160 7.250 4.320 ;
        RECT  7.090 3.060 7.250 4.500 ;
        RECT  6.780 4.160 7.250 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.830 3.790 7.990 4.500 ;
        RECT  6.780 4.340 7.990 4.500 ;
        RECT  7.850 0.560 8.050 2.050 ;
        RECT  7.660 1.440 8.050 2.050 ;
        RECT  7.660 1.770 8.960 2.050 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 9.200 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 9.200 3.660 ;
        RECT  4.820 1.180 9.200 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 9.200 4.800 ;
        RECT  0.000 0.000 9.200 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 9.200 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMQM1HM

MACRO SDFMM8HM
    CLASS CORE ;
    FOREIGN SDFMM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.706  LAYER ME1  ;
        ANTENNADIFFAREA 1.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.770 0.400 9.100 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.071  LAYER ME1  ;
        ANTENNADIFFAREA 1.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.960 4.140 10.300 4.420 ;
        RECT  10.090 2.890 10.300 4.420 ;
        RECT  9.900 2.890 10.300 3.160 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  10.480 1.590 10.640 3.180 ;
        RECT  10.400 1.590 10.640 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  6.010 2.260 6.290 2.720 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  10.440 -0.140 10.640 0.740 ;
        RECT  9.300 -0.140 9.560 0.750 ;
        RECT  8.280 -0.140 8.480 0.700 ;
        RECT  7.240 -0.140 7.460 0.610 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 10.800 4.940 ;
        RECT  10.480 4.020 10.640 4.940 ;
        RECT  9.300 3.970 9.540 4.940 ;
        RECT  8.300 4.240 8.500 4.940 ;
        RECT  6.020 4.480 6.300 4.940 ;
        RECT  3.630 4.320 3.830 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.880 0.320 3.240 ;
        RECT  0.100 2.880 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.130 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.290 ;
        RECT  6.750 3.770 7.100 4.000 ;
        RECT  4.750 3.840 7.100 4.000 ;
        RECT  3.050 4.000 4.230 4.160 ;
        RECT  3.050 4.000 3.390 4.290 ;
        RECT  4.070 4.000 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.810 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.600 2.700 7.810 4.150 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.420 3.360 ;
        RECT  4.850 3.200 7.420 3.360 ;
        RECT  8.430 3.580 8.650 4.080 ;
        RECT  7.970 3.920 8.650 4.080 ;
        RECT  5.070 4.160 7.420 4.320 ;
        RECT  7.260 3.060 7.420 4.500 ;
        RECT  7.010 4.160 7.420 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.970 3.920 8.130 4.500 ;
        RECT  7.010 4.340 8.130 4.500 ;
        RECT  8.750 3.140 9.050 3.360 ;
        RECT  8.810 3.140 9.050 4.470 ;
        RECT  8.010 2.820 9.420 2.980 ;
        RECT  9.240 2.820 9.420 3.810 ;
        RECT  8.010 2.820 8.210 3.630 ;
        RECT  9.240 3.560 9.730 3.810 ;
        RECT  9.310 0.990 9.830 1.240 ;
        RECT  7.780 0.560 7.980 2.060 ;
        RECT  7.660 1.690 7.980 2.060 ;
        RECT  9.310 0.990 9.470 2.060 ;
        RECT  7.660 1.900 9.470 2.060 ;
        RECT  9.900 0.330 10.190 0.830 ;
        RECT  10.010 0.330 10.190 1.990 ;
        RECT  9.900 1.450 10.190 1.990 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 10.800 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 10.800 3.660 ;
        RECT  4.820 1.180 10.800 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 10.800 4.800 ;
        RECT  0.000 0.000 10.800 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 10.800 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMM8HM

MACRO SDFMM4HM
    CLASS CORE ;
    FOREIGN SDFMM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.738  LAYER ME1  ;
        ANTENNADIFFAREA 0.896  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.780 0.550 9.160 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.071  LAYER ME1  ;
        ANTENNADIFFAREA 1.002  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.800 4.140 10.300 4.420 ;
        RECT  10.070 2.900 10.300 4.420 ;
        RECT  9.800 2.900 10.300 3.160 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  6.010 2.260 6.290 2.720 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.330 -0.140 9.490 0.720 ;
        RECT  8.290 -0.140 8.490 0.710 ;
        RECT  7.270 -0.140 7.490 0.440 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 10.400 4.940 ;
        RECT  9.270 4.130 9.530 4.940 ;
        RECT  8.310 4.240 8.510 4.940 ;
        RECT  6.020 4.480 6.300 4.940 ;
        RECT  3.610 4.480 3.890 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.950 0.320 3.300 ;
        RECT  0.100 2.950 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.240 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.250 ;
        RECT  6.750 3.770 7.100 4.000 ;
        RECT  4.750 3.840 7.100 4.000 ;
        RECT  3.050 3.970 4.230 4.250 ;
        RECT  4.070 3.970 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.810 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.600 2.700 7.810 4.150 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.420 3.360 ;
        RECT  4.850 3.200 7.420 3.360 ;
        RECT  8.430 3.580 8.660 4.080 ;
        RECT  7.970 3.920 8.660 4.080 ;
        RECT  5.070 4.160 7.420 4.320 ;
        RECT  7.260 3.060 7.420 4.500 ;
        RECT  7.010 4.160 7.420 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.970 3.920 8.130 4.500 ;
        RECT  7.010 4.340 8.130 4.500 ;
        RECT  8.760 3.140 9.060 3.360 ;
        RECT  8.820 3.140 9.060 4.260 ;
        RECT  8.010 2.820 9.510 2.980 ;
        RECT  9.330 2.820 9.510 3.810 ;
        RECT  8.010 2.820 8.210 3.630 ;
        RECT  9.330 3.560 9.630 3.810 ;
        RECT  9.400 0.980 9.730 1.260 ;
        RECT  7.780 0.560 7.980 2.060 ;
        RECT  7.660 1.480 7.980 2.060 ;
        RECT  9.400 0.980 9.580 2.060 ;
        RECT  7.660 1.900 9.580 2.060 ;
        RECT  9.800 0.330 10.090 0.600 ;
        RECT  9.910 0.330 10.090 1.990 ;
        RECT  9.800 1.700 10.090 1.990 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 10.400 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 10.400 3.660 ;
        RECT  4.820 1.180 10.400 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 10.400 4.800 ;
        RECT  0.000 0.000 10.400 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 10.400 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMM4HM

MACRO SDFMM2HM
    CLASS CORE ;
    FOREIGN SDFMM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.371  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.760 3.080 9.100 3.960 ;
        RECT  8.570 4.130 8.920 4.370 ;
        RECT  8.760 3.080 8.920 4.370 ;
        RECT  8.640 3.080 9.100 3.360 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.411  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.640 4.090 9.900 4.450 ;
        RECT  9.700 2.900 9.900 4.450 ;
        RECT  9.620 2.900 9.900 3.160 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  8.440 -0.140 8.650 0.870 ;
        RECT  7.270 -0.140 7.490 0.440 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 10.000 4.940 ;
        RECT  9.150 4.200 9.310 4.940 ;
        RECT  8.150 4.240 8.350 4.940 ;
        RECT  5.900 4.480 6.180 4.940 ;
        RECT  3.610 4.480 3.890 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.950 0.320 3.300 ;
        RECT  0.100 2.950 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.240 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.250 ;
        RECT  4.750 3.840 6.930 4.000 ;
        RECT  3.050 3.970 4.230 4.250 ;
        RECT  4.070 3.970 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.610 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.410 2.700 7.610 4.160 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.250 3.360 ;
        RECT  4.850 3.200 7.250 3.360 ;
        RECT  8.360 3.580 8.580 3.950 ;
        RECT  7.830 3.790 8.580 3.950 ;
        RECT  5.070 4.160 7.250 4.320 ;
        RECT  7.090 3.060 7.250 4.500 ;
        RECT  6.780 4.160 7.250 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.830 3.790 7.990 4.500 ;
        RECT  6.780 4.340 7.990 4.500 ;
        RECT  7.850 0.560 8.050 2.020 ;
        RECT  7.660 1.540 8.050 2.020 ;
        RECT  7.660 1.860 9.450 2.020 ;
        RECT  7.860 2.700 9.450 2.860 ;
        RECT  9.290 2.700 9.450 3.830 ;
        RECT  7.860 2.700 8.060 3.630 ;
        RECT  9.290 3.550 9.490 3.830 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 10.000 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 10.000 3.660 ;
        RECT  4.820 1.180 10.000 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 10.000 4.800 ;
        RECT  0.000 0.000 10.000 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 10.000 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMM2HM

MACRO SDFMM1HM
    CLASS CORE ;
    FOREIGN SDFMM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.900  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.153  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.450 3.580 1.650 3.780 ;
        LAYER ME2 ;
        RECT  1.300 3.300 1.650 3.960 ;
        LAYER ME1 ;
        RECT  1.380 3.460 1.730 3.920 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 3.500 0.760 3.970 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.940 3.930 1.100 ;
        RECT  1.220 0.900 1.570 1.100 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.950 4.840 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.760 3.080 9.100 3.960 ;
        RECT  8.570 4.260 8.920 4.500 ;
        RECT  8.760 3.080 8.920 4.500 ;
        RECT  8.640 3.080 9.100 3.360 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.640 4.160 9.900 4.500 ;
        RECT  9.700 2.900 9.900 4.500 ;
        RECT  9.620 2.900 9.900 3.160 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 3.480 2.360 3.940 ;
        END
    END S
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.350 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  7.340 1.490 7.500 2.540 ;
        RECT  6.730 1.490 7.500 1.680 ;
        RECT  1.660 2.260 1.880 3.300 ;
        RECT  0.500 3.020 0.840 3.300 ;
        RECT  0.500 2.260 0.660 3.300 ;
        RECT  0.100 1.620 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  8.440 -0.140 8.650 0.870 ;
        RECT  7.270 -0.140 7.490 0.440 ;
        RECT  1.550 -0.140 1.830 0.320 ;
        RECT  0.100 -0.140 0.380 0.660 ;
        RECT  0.000 4.660 10.000 4.940 ;
        RECT  9.150 4.200 9.310 4.940 ;
        RECT  8.150 4.240 8.350 4.940 ;
        RECT  5.900 4.480 6.180 4.940 ;
        RECT  3.610 4.480 3.890 4.940 ;
        RECT  1.930 4.420 2.150 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 2.700 1.190 2.860 ;
        RECT  1.000 2.700 1.190 4.180 ;
        RECT  1.000 3.020 1.330 3.300 ;
        RECT  1.000 3.020 1.210 4.180 ;
        RECT  0.760 0.850 0.980 1.460 ;
        RECT  0.760 1.300 1.880 1.460 ;
        RECT  0.100 2.950 0.320 3.300 ;
        RECT  0.100 2.950 0.260 4.500 ;
        RECT  1.590 4.100 2.470 4.260 ;
        RECT  0.100 4.240 0.410 4.500 ;
        RECT  2.310 4.100 2.470 4.500 ;
        RECT  1.590 4.100 1.750 4.500 ;
        RECT  0.100 4.340 1.750 4.500 ;
        RECT  2.310 4.340 2.830 4.500 ;
        RECT  2.310 2.700 2.620 3.300 ;
        RECT  2.240 3.020 2.620 3.300 ;
        RECT  2.240 3.140 2.830 3.300 ;
        RECT  2.630 3.140 2.830 4.180 ;
        RECT  1.830 1.620 4.300 1.780 ;
        RECT  4.100 0.950 4.320 1.460 ;
        RECT  2.270 1.300 4.320 1.460 ;
        RECT  2.330 0.620 5.120 0.780 ;
        RECT  0.940 1.620 1.220 2.100 ;
        RECT  0.940 1.940 5.440 2.100 ;
        RECT  1.990 0.300 5.560 0.460 ;
        RECT  5.260 0.300 5.560 0.530 ;
        RECT  1.990 0.300 2.160 0.660 ;
        RECT  0.890 0.500 2.160 0.660 ;
        RECT  4.340 3.020 4.650 3.280 ;
        RECT  4.390 3.020 4.650 3.680 ;
        RECT  4.390 3.520 6.110 3.680 ;
        RECT  4.390 3.020 4.590 4.180 ;
        RECT  5.800 0.310 6.080 0.870 ;
        RECT  5.280 0.710 6.080 0.870 ;
        RECT  5.280 0.710 5.440 1.660 ;
        RECT  5.120 1.320 5.440 1.660 ;
        RECT  5.120 1.500 6.160 1.660 ;
        RECT  3.050 3.000 3.410 3.280 ;
        RECT  3.050 3.000 3.230 4.250 ;
        RECT  4.750 3.840 6.930 4.000 ;
        RECT  3.050 3.970 4.230 4.250 ;
        RECT  4.070 3.970 4.230 4.500 ;
        RECT  4.750 3.840 4.910 4.500 ;
        RECT  4.070 4.340 4.910 4.500 ;
        RECT  6.020 1.860 7.180 2.060 ;
        RECT  6.590 0.710 6.790 1.270 ;
        RECT  6.590 1.060 7.600 1.270 ;
        RECT  7.340 0.990 7.600 1.270 ;
        RECT  5.600 1.110 7.600 1.270 ;
        RECT  3.570 2.700 5.580 2.860 ;
        RECT  6.480 2.700 7.610 2.860 ;
        RECT  5.420 2.700 5.580 3.040 ;
        RECT  6.480 2.700 6.640 3.040 ;
        RECT  5.420 2.880 6.640 3.040 ;
        RECT  3.570 2.700 3.730 3.790 ;
        RECT  3.390 3.500 3.730 3.790 ;
        RECT  7.410 2.700 7.610 4.160 ;
        RECT  4.850 3.060 5.130 3.360 ;
        RECT  6.880 3.060 7.250 3.360 ;
        RECT  4.850 3.200 7.250 3.360 ;
        RECT  8.360 3.580 8.580 3.950 ;
        RECT  7.830 3.790 8.580 3.950 ;
        RECT  5.070 4.160 7.250 4.320 ;
        RECT  7.090 3.060 7.250 4.500 ;
        RECT  6.780 4.160 7.250 4.500 ;
        RECT  5.070 4.160 5.270 4.470 ;
        RECT  7.830 3.790 7.990 4.500 ;
        RECT  6.780 4.340 7.990 4.500 ;
        RECT  7.850 0.560 8.050 2.020 ;
        RECT  7.660 1.540 8.050 2.020 ;
        RECT  7.660 1.860 9.450 2.020 ;
        RECT  7.860 2.700 9.450 2.860 ;
        RECT  9.290 2.700 9.450 3.830 ;
        RECT  7.860 2.700 8.060 3.630 ;
        RECT  9.290 3.550 9.490 3.830 ;
        LAYER VTPH ;
        RECT  5.250 1.100 7.330 3.660 ;
        RECT  0.000 1.140 0.930 3.600 ;
        RECT  0.000 1.180 10.000 3.580 ;
        RECT  0.000 1.180 2.940 3.600 ;
        RECT  0.000 1.140 0.770 3.660 ;
        RECT  5.250 1.140 10.000 3.660 ;
        RECT  4.820 1.180 10.000 3.660 ;
        LAYER VTNH ;
        RECT  2.940 3.580 4.820 4.800 ;
        RECT  0.770 3.600 4.820 4.800 ;
        RECT  0.000 3.660 10.000 4.800 ;
        RECT  0.000 0.000 10.000 1.100 ;
        RECT  0.000 0.000 5.250 1.140 ;
        RECT  7.330 0.000 10.000 1.140 ;
        RECT  0.930 0.000 5.250 1.180 ;
    END
END SDFMM1HM

MACRO SDFM8HM
    CLASS CORE ;
    FOREIGN SDFM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.884  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.900 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.010 1.200 1.380 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.214  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.330 1.100 3.530 1.300 ;
        LAYER ME2 ;
        RECT  3.300 0.900 3.560 1.560 ;
        LAYER ME1 ;
        RECT  3.220 1.060 3.850 1.320 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.744  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.480 1.100 2.680 1.300 ;
        LAYER ME2 ;
        RECT  2.450 0.900 2.710 1.560 ;
        LAYER ME1 ;
        RECT  2.320 0.980 2.680 1.380 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.068  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.550 0.800 14.350 0.960 ;
        RECT  14.070 0.620 14.350 0.960 ;
        RECT  13.600 0.800 13.900 1.680 ;
        RECT  12.550 0.620 12.830 1.680 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.890 0.390 18.090 2.100 ;
        RECT  16.840 0.840 18.090 1.100 ;
        RECT  16.840 0.390 17.070 2.100 ;
        END
    END QB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.188  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.360 0.660 1.560 0.970 ;
        RECT  0.500 0.660 1.560 0.850 ;
        RECT  0.500 0.660 0.700 1.190 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.800 2.540 ;
        RECT  18.410 1.460 18.610 2.540 ;
        RECT  17.370 1.460 17.570 2.540 ;
        RECT  16.270 1.470 16.470 2.540 ;
        RECT  14.410 2.080 14.690 2.540 ;
        RECT  8.110 1.860 8.390 2.540 ;
        RECT  4.860 1.970 5.020 2.540 ;
        RECT  3.480 1.800 3.680 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.800 0.140 ;
        RECT  18.420 -0.140 18.620 0.670 ;
        RECT  17.370 -0.140 17.570 0.670 ;
        RECT  16.350 -0.140 16.510 0.710 ;
        RECT  14.830 -0.140 15.110 0.320 ;
        RECT  13.310 -0.140 13.590 0.320 ;
        RECT  11.870 -0.140 12.070 0.380 ;
        RECT  10.910 -0.140 11.190 0.560 ;
        RECT  7.920 -0.140 8.200 0.340 ;
        RECT  4.940 -0.140 5.100 0.420 ;
        RECT  3.480 -0.140 3.680 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.820 0.820 2.020 1.700 ;
        RECT  0.140 1.540 2.020 1.700 ;
        RECT  0.140 0.300 0.340 2.100 ;
        RECT  2.210 0.620 3.000 0.820 ;
        RECT  2.840 0.620 3.000 1.700 ;
        RECT  2.260 1.540 3.000 1.700 ;
        RECT  4.160 0.620 4.440 1.200 ;
        RECT  4.160 1.000 5.230 1.200 ;
        RECT  4.160 0.620 4.380 1.760 ;
        RECT  5.580 0.620 5.860 1.540 ;
        RECT  5.500 1.340 6.310 1.540 ;
        RECT  5.500 1.340 5.770 1.780 ;
        RECT  3.160 1.480 4.000 1.640 ;
        RECT  4.540 1.550 5.340 1.710 ;
        RECT  3.840 1.480 4.000 2.100 ;
        RECT  5.180 1.550 5.340 2.100 ;
        RECT  3.160 1.480 3.320 2.020 ;
        RECT  1.550 1.860 3.320 2.020 ;
        RECT  4.540 1.550 4.700 2.100 ;
        RECT  3.840 1.940 4.700 2.100 ;
        RECT  6.040 1.900 6.320 2.100 ;
        RECT  5.180 1.940 6.320 2.100 ;
        RECT  1.550 0.300 3.320 0.460 ;
        RECT  3.840 0.300 4.760 0.460 ;
        RECT  5.260 0.300 6.450 0.460 ;
        RECT  1.550 0.300 1.830 0.500 ;
        RECT  6.090 0.300 6.450 0.560 ;
        RECT  4.600 0.300 4.760 0.740 ;
        RECT  3.160 0.300 3.320 0.880 ;
        RECT  5.260 0.300 5.420 0.740 ;
        RECT  4.600 0.580 5.420 0.740 ;
        RECT  3.840 0.300 4.000 0.880 ;
        RECT  3.160 0.720 4.000 0.880 ;
        RECT  6.090 0.820 6.640 1.100 ;
        RECT  6.480 0.820 6.640 2.100 ;
        RECT  7.260 1.480 7.480 2.100 ;
        RECT  6.480 1.940 7.480 2.100 ;
        RECT  6.670 0.300 6.960 0.570 ;
        RECT  7.560 0.840 8.350 1.000 ;
        RECT  6.800 0.300 6.960 1.780 ;
        RECT  7.560 0.840 7.720 1.200 ;
        RECT  6.800 1.040 7.720 1.200 ;
        RECT  6.800 1.040 7.050 1.780 ;
        RECT  7.890 1.280 9.140 1.480 ;
        RECT  8.860 0.620 9.140 1.750 ;
        RECT  8.750 1.280 9.140 1.750 ;
        RECT  8.380 0.300 10.150 0.460 ;
        RECT  8.380 0.300 8.540 0.660 ;
        RECT  7.120 0.500 8.540 0.660 ;
        RECT  7.120 0.500 7.400 0.880 ;
        RECT  9.990 0.300 10.150 1.780 ;
        RECT  9.930 1.560 10.210 1.780 ;
        RECT  9.450 0.620 9.830 0.900 ;
        RECT  15.150 1.120 15.430 1.920 ;
        RECT  14.090 1.760 15.430 1.920 ;
        RECT  9.450 0.620 9.610 2.100 ;
        RECT  14.090 1.760 14.250 2.100 ;
        RECT  9.450 1.940 14.250 2.100 ;
        RECT  15.590 0.620 15.870 0.960 ;
        RECT  14.510 0.800 15.870 0.960 ;
        RECT  14.510 0.800 14.670 1.320 ;
        RECT  14.130 1.120 14.670 1.320 ;
        RECT  15.650 0.620 15.870 2.100 ;
        RECT  12.230 0.300 13.150 0.460 ;
        RECT  13.750 0.300 14.670 0.460 ;
        RECT  15.270 0.300 16.190 0.460 ;
        RECT  12.990 0.300 13.150 0.640 ;
        RECT  14.510 0.300 14.670 0.640 ;
        RECT  13.750 0.300 13.910 0.640 ;
        RECT  12.990 0.480 13.910 0.640 ;
        RECT  15.270 0.300 15.430 0.640 ;
        RECT  14.510 0.480 15.430 0.640 ;
        RECT  10.370 0.410 10.570 1.660 ;
        RECT  11.470 0.540 11.670 0.880 ;
        RECT  12.230 0.300 12.390 0.880 ;
        RECT  10.370 0.720 12.390 0.880 ;
        RECT  16.030 0.300 16.190 1.230 ;
        RECT  16.030 1.030 16.670 1.230 ;
        RECT  10.370 0.720 10.670 1.660 ;
        RECT  10.370 1.500 11.700 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.460 2.400 ;
        RECT  10.040 1.140 18.800 2.400 ;
        RECT  0.000 1.200 18.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.800 1.140 ;
        RECT  8.460 0.000 10.040 1.200 ;
    END
END SDFM8HM

MACRO SDFM4HM
    CLASS CORE ;
    FOREIGN SDFM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.884  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.900 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.010 1.200 1.380 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.026  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.330 1.100 3.530 1.300 ;
        LAYER ME2 ;
        RECT  3.300 0.900 3.560 1.560 ;
        LAYER ME1 ;
        RECT  3.220 1.060 3.850 1.320 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.656  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.480 1.100 2.680 1.300 ;
        LAYER ME2 ;
        RECT  2.450 0.900 2.710 1.560 ;
        LAYER ME1 ;
        RECT  2.320 0.980 2.680 1.380 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.648  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.240 1.240 11.830 1.680 ;
        RECT  11.550 0.620 11.830 1.680 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.320 0.390 14.700 2.100 ;
        END
    END QB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.186  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.360 0.660 1.560 0.970 ;
        RECT  0.500 0.660 1.560 0.850 ;
        RECT  0.500 0.660 0.700 1.190 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.870 1.820 15.070 2.540 ;
        RECT  13.750 1.470 13.950 2.540 ;
        RECT  12.410 2.020 12.630 2.540 ;
        RECT  8.110 1.860 8.390 2.540 ;
        RECT  4.860 1.970 5.020 2.540 ;
        RECT  3.480 1.800 3.680 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.870 -0.140 15.070 0.670 ;
        RECT  13.830 -0.140 13.990 0.710 ;
        RECT  12.310 -0.140 12.590 0.320 ;
        RECT  10.850 -0.140 11.070 0.640 ;
        RECT  7.920 -0.140 8.200 0.340 ;
        RECT  4.940 -0.140 5.100 0.420 ;
        RECT  3.480 -0.140 3.680 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.350 0.380 0.550 ;
        RECT  0.100 0.350 0.330 2.100 ;
        RECT  1.820 0.820 2.020 1.700 ;
        RECT  0.100 1.540 2.020 1.700 ;
        RECT  0.100 1.540 0.340 2.100 ;
        RECT  2.210 0.620 3.000 0.820 ;
        RECT  2.840 0.620 3.000 1.700 ;
        RECT  2.260 1.540 3.000 1.700 ;
        RECT  4.160 0.620 4.440 1.200 ;
        RECT  4.160 1.000 5.230 1.200 ;
        RECT  4.160 0.620 4.380 1.760 ;
        RECT  5.580 0.620 5.860 1.540 ;
        RECT  5.500 1.340 6.310 1.540 ;
        RECT  5.500 1.340 5.770 1.780 ;
        RECT  3.160 1.480 4.000 1.640 ;
        RECT  4.540 1.550 5.340 1.710 ;
        RECT  3.840 1.480 4.000 2.100 ;
        RECT  5.180 1.550 5.340 2.100 ;
        RECT  3.160 1.480 3.320 2.020 ;
        RECT  1.550 1.860 3.320 2.020 ;
        RECT  4.540 1.550 4.700 2.100 ;
        RECT  3.840 1.940 4.700 2.100 ;
        RECT  6.040 1.900 6.320 2.100 ;
        RECT  5.180 1.940 6.320 2.100 ;
        RECT  1.550 0.300 3.320 0.460 ;
        RECT  3.840 0.300 4.760 0.460 ;
        RECT  5.260 0.300 6.450 0.460 ;
        RECT  1.550 0.300 1.830 0.500 ;
        RECT  6.090 0.300 6.450 0.560 ;
        RECT  4.600 0.300 4.760 0.740 ;
        RECT  3.160 0.300 3.320 0.880 ;
        RECT  5.260 0.300 5.420 0.740 ;
        RECT  4.600 0.580 5.420 0.740 ;
        RECT  3.840 0.300 4.000 0.880 ;
        RECT  3.160 0.720 4.000 0.880 ;
        RECT  6.090 0.820 6.640 1.100 ;
        RECT  6.480 0.820 6.640 2.100 ;
        RECT  7.260 1.480 7.480 2.100 ;
        RECT  6.480 1.940 7.480 2.100 ;
        RECT  6.670 0.300 6.960 0.570 ;
        RECT  7.560 0.840 8.350 1.000 ;
        RECT  6.800 0.300 6.960 1.780 ;
        RECT  7.560 0.840 7.720 1.200 ;
        RECT  6.800 1.040 7.720 1.200 ;
        RECT  6.800 1.040 7.050 1.780 ;
        RECT  7.890 1.280 9.140 1.480 ;
        RECT  8.860 0.620 9.140 1.750 ;
        RECT  8.750 1.280 9.140 1.750 ;
        RECT  8.380 0.300 10.210 0.460 ;
        RECT  8.380 0.300 8.540 0.660 ;
        RECT  7.120 0.500 8.540 0.660 ;
        RECT  7.120 0.500 7.400 0.880 ;
        RECT  9.990 0.300 10.210 1.780 ;
        RECT  9.930 1.560 10.210 1.780 ;
        RECT  9.450 0.620 9.830 0.900 ;
        RECT  12.530 1.120 12.810 1.780 ;
        RECT  12.090 1.620 12.810 1.780 ;
        RECT  9.450 0.620 9.610 2.100 ;
        RECT  12.090 1.620 12.250 2.100 ;
        RECT  9.450 1.940 12.250 2.100 ;
        RECT  13.070 0.620 13.350 0.960 ;
        RECT  11.990 0.800 13.350 0.960 ;
        RECT  11.990 0.800 12.190 1.280 ;
        RECT  13.130 0.620 13.350 2.100 ;
        RECT  11.230 0.300 12.150 0.460 ;
        RECT  12.750 0.300 13.670 0.460 ;
        RECT  11.990 0.300 12.150 0.640 ;
        RECT  12.750 0.300 12.910 0.640 ;
        RECT  11.990 0.480 12.910 0.640 ;
        RECT  10.370 0.410 10.600 1.720 ;
        RECT  11.230 0.300 11.390 1.000 ;
        RECT  10.370 0.840 11.390 1.000 ;
        RECT  13.510 0.300 13.670 1.230 ;
        RECT  13.510 1.030 14.150 1.230 ;
        RECT  10.370 0.840 10.610 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.460 2.400 ;
        RECT  10.040 1.140 15.200 2.400 ;
        RECT  0.000 1.200 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 1.140 ;
        RECT  8.460 0.000 10.040 1.200 ;
    END
END SDFM4HM

MACRO SDFM2HM
    CLASS CORE ;
    FOREIGN SDFM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.884  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.900 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.010 1.200 1.380 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.026  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.330 1.100 3.530 1.300 ;
        LAYER ME2 ;
        RECT  3.300 0.900 3.560 1.560 ;
        LAYER ME1 ;
        RECT  3.220 1.060 3.850 1.320 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.656  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.480 1.100 2.680 1.300 ;
        LAYER ME2 ;
        RECT  2.450 0.900 2.710 1.560 ;
        LAYER ME1 ;
        RECT  2.320 0.980 2.680 1.380 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.434  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.840 1.240 11.550 1.400 ;
        RECT  11.270 0.620 11.550 1.400 ;
        RECT  10.840 1.240 11.250 1.760 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.427  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.560 0.390 13.900 2.100 ;
        END
    END QB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.186  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.360 0.660 1.560 0.970 ;
        RECT  0.500 0.660 1.560 0.850 ;
        RECT  0.500 0.660 0.700 1.190 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.010 1.470 13.210 2.540 ;
        RECT  11.730 1.980 11.890 2.540 ;
        RECT  8.040 1.860 8.320 2.540 ;
        RECT  4.860 1.970 5.020 2.540 ;
        RECT  3.480 1.800 3.680 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.070 -0.140 13.230 0.710 ;
        RECT  10.570 -0.140 10.790 0.640 ;
        RECT  7.850 -0.140 8.130 0.340 ;
        RECT  4.940 -0.140 5.100 0.420 ;
        RECT  3.480 -0.140 3.680 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.350 0.380 0.550 ;
        RECT  0.100 0.350 0.330 2.100 ;
        RECT  1.820 0.820 2.020 1.700 ;
        RECT  0.100 1.540 2.020 1.700 ;
        RECT  0.100 1.540 0.340 2.100 ;
        RECT  2.210 0.620 3.000 0.820 ;
        RECT  2.840 0.620 3.000 1.700 ;
        RECT  2.260 1.540 3.000 1.700 ;
        RECT  4.160 0.620 4.440 1.200 ;
        RECT  4.160 1.000 5.230 1.200 ;
        RECT  4.160 0.620 4.380 1.760 ;
        RECT  5.580 0.620 5.860 1.540 ;
        RECT  5.500 1.340 6.240 1.540 ;
        RECT  5.500 1.340 5.770 1.780 ;
        RECT  3.160 1.480 4.000 1.640 ;
        RECT  4.540 1.550 5.340 1.710 ;
        RECT  3.840 1.480 4.000 2.100 ;
        RECT  5.180 1.550 5.340 2.100 ;
        RECT  3.160 1.480 3.320 2.020 ;
        RECT  1.550 1.860 3.320 2.020 ;
        RECT  4.540 1.550 4.700 2.100 ;
        RECT  3.840 1.940 4.700 2.100 ;
        RECT  5.970 1.900 6.250 2.100 ;
        RECT  5.180 1.940 6.250 2.100 ;
        RECT  1.550 0.300 3.320 0.460 ;
        RECT  3.840 0.300 4.760 0.460 ;
        RECT  5.260 0.300 6.380 0.460 ;
        RECT  1.550 0.300 1.830 0.500 ;
        RECT  6.020 0.300 6.380 0.560 ;
        RECT  4.600 0.300 4.760 0.740 ;
        RECT  3.160 0.300 3.320 0.880 ;
        RECT  5.260 0.300 5.420 0.740 ;
        RECT  4.600 0.580 5.420 0.740 ;
        RECT  3.840 0.300 4.000 0.880 ;
        RECT  3.160 0.720 4.000 0.880 ;
        RECT  6.020 0.820 6.570 1.100 ;
        RECT  6.410 0.820 6.570 2.100 ;
        RECT  7.190 1.480 7.410 2.100 ;
        RECT  6.410 1.940 7.410 2.100 ;
        RECT  6.600 0.300 6.890 0.570 ;
        RECT  7.490 0.840 8.280 1.000 ;
        RECT  6.730 0.300 6.890 1.780 ;
        RECT  7.490 0.840 7.650 1.200 ;
        RECT  6.730 1.040 7.650 1.200 ;
        RECT  6.730 1.040 6.980 1.780 ;
        RECT  7.820 1.280 9.070 1.480 ;
        RECT  8.790 0.620 9.070 1.750 ;
        RECT  8.660 1.280 9.070 1.750 ;
        RECT  8.310 0.300 9.930 0.460 ;
        RECT  8.310 0.300 8.470 0.660 ;
        RECT  7.050 0.500 8.470 0.660 ;
        RECT  7.050 0.500 7.330 0.880 ;
        RECT  9.690 0.300 9.930 1.780 ;
        RECT  9.650 1.560 9.930 1.780 ;
        RECT  9.240 0.620 9.530 0.900 ;
        RECT  11.410 1.620 11.790 1.780 ;
        RECT  9.240 0.620 9.400 2.100 ;
        RECT  11.410 1.620 11.570 2.100 ;
        RECT  9.240 1.940 11.570 2.100 ;
        RECT  12.050 0.560 12.650 0.840 ;
        RECT  12.370 0.560 12.530 1.760 ;
        RECT  10.950 0.300 11.870 0.460 ;
        RECT  10.090 0.300 10.320 1.720 ;
        RECT  10.950 0.300 11.110 1.000 ;
        RECT  10.090 0.840 11.110 1.000 ;
        RECT  12.690 1.030 13.390 1.230 ;
        RECT  11.710 0.300 11.870 1.400 ;
        RECT  11.710 1.240 12.210 1.400 ;
        RECT  10.090 0.840 10.330 1.720 ;
        RECT  12.050 1.240 12.210 2.100 ;
        RECT  12.690 1.030 12.850 2.100 ;
        RECT  12.050 1.940 12.850 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.390 2.400 ;
        RECT  9.830 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.140 ;
        RECT  8.390 0.000 9.830 1.200 ;
    END
END SDFM2HM

MACRO SDFM1HM
    CLASS CORE ;
    FOREIGN SDFM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.884  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.930 1.100 1.130 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.010 1.200 1.380 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        ANTENNAGATEAREA 0.056  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.206  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.000 1.100 3.200 1.300 ;
        LAYER ME2 ;
        RECT  2.900 0.900 3.200 1.560 ;
        LAYER ME1 ;
        RECT  2.890 1.060 3.520 1.320 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.228  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.050 1.100 2.250 1.300 ;
        LAYER ME2 ;
        RECT  2.050 0.900 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.890 0.980 2.250 1.380 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.393  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.440 1.240 11.220 1.400 ;
        RECT  10.940 0.620 11.220 1.400 ;
        RECT  10.440 1.240 10.920 1.760 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.368  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.230 0.300 13.500 2.100 ;
        END
    END QB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.410 0.660 1.610 0.970 ;
        RECT  0.500 0.660 1.610 0.850 ;
        RECT  0.500 0.660 0.700 1.190 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.680 1.470 12.880 2.540 ;
        RECT  11.400 1.980 11.560 2.540 ;
        RECT  7.710 1.860 7.990 2.540 ;
        RECT  4.530 1.970 4.690 2.540 ;
        RECT  3.150 1.800 3.350 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.680 -0.140 12.900 0.620 ;
        RECT  10.240 -0.140 10.460 0.640 ;
        RECT  7.520 -0.140 7.800 0.340 ;
        RECT  4.610 -0.140 4.770 0.420 ;
        RECT  3.150 -0.140 3.350 0.560 ;
        RECT  0.650 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.350 0.380 0.550 ;
        RECT  0.100 0.350 0.330 2.100 ;
        RECT  1.440 1.180 1.640 1.700 ;
        RECT  2.470 0.640 2.670 1.700 ;
        RECT  0.100 1.540 2.670 1.700 ;
        RECT  0.100 1.540 0.340 2.100 ;
        RECT  3.830 0.620 4.110 1.200 ;
        RECT  3.830 1.000 4.900 1.200 ;
        RECT  3.830 0.620 4.050 1.760 ;
        RECT  5.250 0.620 5.530 1.540 ;
        RECT  5.170 1.340 5.910 1.540 ;
        RECT  5.170 1.340 5.440 1.780 ;
        RECT  2.830 1.480 3.670 1.640 ;
        RECT  4.210 1.550 5.010 1.710 ;
        RECT  3.510 1.480 3.670 2.100 ;
        RECT  4.850 1.550 5.010 2.100 ;
        RECT  2.830 1.480 2.990 2.020 ;
        RECT  1.600 1.860 2.990 2.020 ;
        RECT  4.210 1.550 4.370 2.100 ;
        RECT  3.510 1.940 4.370 2.100 ;
        RECT  5.640 1.900 5.920 2.100 ;
        RECT  4.850 1.940 5.920 2.100 ;
        RECT  1.700 0.300 2.990 0.460 ;
        RECT  3.510 0.300 4.430 0.460 ;
        RECT  4.930 0.300 6.050 0.460 ;
        RECT  1.700 0.300 1.980 0.500 ;
        RECT  5.690 0.300 6.050 0.560 ;
        RECT  4.270 0.300 4.430 0.740 ;
        RECT  2.830 0.300 2.990 0.880 ;
        RECT  4.930 0.300 5.090 0.740 ;
        RECT  4.270 0.580 5.090 0.740 ;
        RECT  3.510 0.300 3.670 0.880 ;
        RECT  2.830 0.720 3.670 0.880 ;
        RECT  5.690 0.820 6.240 1.100 ;
        RECT  6.080 0.820 6.240 2.100 ;
        RECT  6.860 1.480 7.080 2.100 ;
        RECT  6.080 1.940 7.080 2.100 ;
        RECT  6.270 0.300 6.560 0.570 ;
        RECT  7.160 0.840 7.950 1.000 ;
        RECT  6.400 0.300 6.560 1.780 ;
        RECT  7.160 0.840 7.320 1.200 ;
        RECT  6.400 1.040 7.320 1.200 ;
        RECT  6.400 1.040 6.650 1.780 ;
        RECT  7.490 1.280 8.740 1.480 ;
        RECT  8.460 0.620 8.740 1.750 ;
        RECT  8.330 1.280 8.740 1.750 ;
        RECT  7.980 0.300 9.520 0.460 ;
        RECT  7.980 0.300 8.140 0.660 ;
        RECT  6.720 0.500 8.140 0.660 ;
        RECT  6.720 0.500 7.000 0.880 ;
        RECT  9.360 0.300 9.520 1.780 ;
        RECT  9.320 1.560 9.600 1.780 ;
        RECT  8.910 0.620 9.200 0.900 ;
        RECT  11.080 1.620 11.460 1.780 ;
        RECT  8.910 0.620 9.070 2.100 ;
        RECT  11.080 1.620 11.240 2.100 ;
        RECT  8.910 1.940 11.240 2.100 ;
        RECT  11.720 0.300 12.320 0.570 ;
        RECT  11.720 0.300 12.200 0.580 ;
        RECT  12.040 0.300 12.200 1.760 ;
        RECT  10.620 0.300 11.540 0.460 ;
        RECT  9.680 0.300 9.990 0.660 ;
        RECT  9.760 0.300 9.990 1.720 ;
        RECT  10.620 0.300 10.780 1.000 ;
        RECT  9.760 0.840 10.780 1.000 ;
        RECT  12.360 1.030 13.060 1.230 ;
        RECT  11.380 0.300 11.540 1.400 ;
        RECT  11.380 1.240 11.880 1.400 ;
        RECT  9.760 0.840 10.000 1.720 ;
        RECT  11.720 1.240 11.880 2.100 ;
        RECT  12.360 1.030 12.520 2.100 ;
        RECT  11.720 1.940 12.520 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.060 2.400 ;
        RECT  9.500 1.140 13.600 2.400 ;
        RECT  0.000 1.200 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.140 ;
        RECT  8.060 0.000 9.500 1.200 ;
    END
END SDFM1HM

MACRO SDFEZRM8HM
    CLASS CORE ;
    FOREIGN SDFEZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 3.570 3.720 3.900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 0.840 1.900 1.200 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 0.720 1.250 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.794  LAYER ME1  ;
        ANTENNADIFFAREA 1.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.620 3.080 9.900 4.420 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.981  LAYER ME1  ;
        ANTENNADIFFAREA 1.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.700 4.180 11.100 4.380 ;
        RECT  10.900 3.070 11.100 4.380 ;
        RECT  10.700 3.070 11.100 3.270 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.620 0.900 5.160 1.220 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.047  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.110 2.760 1.500 3.160 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 3.640 2.560 3.800 ;
        RECT  2.400 3.420 2.560 3.800 ;
        RECT  0.500 3.920 1.720 4.080 ;
        RECT  1.560 3.640 1.720 4.080 ;
        RECT  0.500 3.640 0.700 4.080 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.260 1.480 11.460 3.340 ;
        RECT  7.900 2.140 8.180 2.540 ;
        RECT  7.940 2.140 8.140 3.340 ;
        RECT  7.400 2.260 7.600 3.430 ;
        RECT  0.660 1.730 0.940 2.540 ;
        RECT  0.700 1.730 0.900 3.160 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.260 -0.140 11.460 0.610 ;
        RECT  10.180 -0.140 10.380 0.610 ;
        RECT  9.060 -0.140 9.260 0.610 ;
        RECT  7.980 -0.140 8.180 0.560 ;
        RECT  7.460 -0.140 7.660 0.560 ;
        RECT  4.460 -0.140 4.660 0.420 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 11.600 4.940 ;
        RECT  11.260 4.240 11.460 4.940 ;
        RECT  10.180 4.240 10.380 4.940 ;
        RECT  9.060 4.240 9.260 4.940 ;
        RECT  7.940 4.240 8.140 4.940 ;
        RECT  7.380 4.240 7.580 4.940 ;
        RECT  5.240 4.240 5.440 4.940 ;
        RECT  3.360 4.380 3.520 4.940 ;
        RECT  0.660 4.480 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.660 2.760 1.860 3.480 ;
        RECT  0.140 3.320 1.860 3.480 ;
        RECT  0.140 3.040 0.340 4.480 ;
        RECT  2.060 0.960 2.800 1.120 ;
        RECT  0.960 0.950 1.160 1.570 ;
        RECT  2.060 0.960 2.220 1.570 ;
        RECT  0.140 1.410 2.220 1.570 ;
        RECT  0.140 0.320 0.340 1.910 ;
        RECT  2.520 3.040 2.880 3.240 ;
        RECT  2.720 3.040 2.880 4.160 ;
        RECT  2.140 4.000 2.880 4.160 ;
        RECT  2.060 0.640 3.120 0.800 ;
        RECT  2.960 1.020 3.560 1.220 ;
        RECT  2.960 0.640 3.120 1.440 ;
        RECT  2.380 1.280 3.120 1.440 ;
        RECT  2.380 1.280 2.540 2.070 ;
        RECT  1.620 1.870 2.540 2.070 ;
        RECT  3.620 0.640 3.980 0.800 ;
        RECT  3.780 0.640 3.980 1.760 ;
        RECT  2.920 1.600 3.980 1.760 ;
        RECT  2.920 1.600 3.120 2.080 ;
        RECT  3.660 3.040 4.280 3.240 ;
        RECT  4.000 3.040 4.280 4.160 ;
        RECT  1.140 0.320 4.300 0.480 ;
        RECT  4.140 0.320 4.300 0.740 ;
        RECT  1.140 0.320 1.340 0.600 ;
        RECT  5.040 0.370 5.200 0.740 ;
        RECT  4.140 0.580 5.200 0.740 ;
        RECT  4.140 0.940 4.300 1.760 ;
        RECT  4.140 1.600 5.300 1.760 ;
        RECT  2.040 2.720 5.660 2.880 ;
        RECT  5.460 2.720 5.660 3.110 ;
        RECT  2.040 2.720 2.240 3.170 ;
        RECT  4.920 3.920 5.920 4.080 ;
        RECT  3.040 4.060 3.840 4.220 ;
        RECT  3.680 4.060 3.840 4.480 ;
        RECT  5.720 3.920 5.920 4.430 ;
        RECT  3.040 4.060 3.200 4.480 ;
        RECT  1.540 4.320 3.200 4.480 ;
        RECT  4.920 3.920 5.080 4.480 ;
        RECT  3.680 4.320 5.080 4.480 ;
        RECT  4.980 3.060 5.180 3.540 ;
        RECT  4.480 3.380 6.620 3.540 ;
        RECT  6.460 3.380 6.620 4.070 ;
        RECT  4.480 3.380 4.760 4.160 ;
        RECT  5.980 2.720 6.940 2.920 ;
        RECT  5.980 2.720 6.180 3.110 ;
        RECT  6.780 2.720 6.940 4.460 ;
        RECT  6.220 4.300 6.940 4.460 ;
        RECT  6.700 1.330 7.720 1.490 ;
        RECT  6.700 0.660 6.980 1.750 ;
        RECT  6.020 0.340 7.300 0.500 ;
        RECT  7.140 0.340 7.300 1.170 ;
        RECT  7.140 0.970 8.440 1.170 ;
        RECT  6.020 0.340 6.180 1.730 ;
        RECT  6.020 1.570 6.500 1.730 ;
        RECT  8.420 0.390 8.780 0.550 ;
        RECT  8.620 0.970 9.400 1.170 ;
        RECT  8.620 0.390 8.780 1.660 ;
        RECT  8.420 1.500 8.780 1.660 ;
        RECT  9.540 0.390 9.900 0.550 ;
        RECT  9.740 0.390 9.900 1.660 ;
        RECT  9.540 1.500 9.900 1.660 ;
        RECT  5.460 0.320 5.820 0.520 ;
        RECT  5.620 0.320 5.820 2.080 ;
        RECT  7.140 1.820 10.580 1.980 ;
        RECT  5.620 1.910 10.580 1.980 ;
        RECT  10.380 0.930 10.580 1.980 ;
        RECT  3.320 1.920 7.300 2.080 ;
        RECT  8.500 2.760 10.310 2.920 ;
        RECT  10.150 2.760 10.310 3.780 ;
        RECT  10.150 3.580 10.590 3.780 ;
        RECT  8.500 2.760 8.700 4.420 ;
        RECT  10.740 0.380 10.940 2.080 ;
        LAYER VTPH ;
        RECT  2.500 1.140 3.300 3.640 ;
        RECT  0.000 1.160 6.400 3.640 ;
        RECT  4.050 1.140 6.400 3.640 ;
        RECT  0.000 1.140 1.850 3.660 ;
        RECT  2.650 1.160 3.750 3.660 ;
        RECT  7.250 1.140 11.600 3.660 ;
        RECT  5.750 1.180 7.820 3.730 ;
        RECT  0.630 1.160 1.900 3.810 ;
        LAYER VTNH ;
        RECT  1.900 3.640 2.650 4.800 ;
        RECT  3.750 3.640 5.750 4.800 ;
        RECT  1.900 3.660 5.750 4.800 ;
        RECT  0.000 3.660 0.630 4.800 ;
        RECT  1.900 3.730 11.600 4.800 ;
        RECT  7.820 3.660 11.600 4.800 ;
        RECT  0.000 3.810 11.600 4.800 ;
        RECT  0.000 0.000 11.600 1.140 ;
        RECT  1.850 0.000 2.500 1.160 ;
        RECT  3.300 0.000 4.050 1.160 ;
        RECT  6.400 0.000 7.250 1.180 ;
    END
END SDFEZRM8HM

MACRO SDFEZRM4HM
    CLASS CORE ;
    FOREIGN SDFEZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 3.570 3.720 3.900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 0.840 1.900 1.210 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 0.720 1.250 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.272  LAYER ME1  ;
        ANTENNADIFFAREA 0.978  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.980 3.980 9.680 4.140 ;
        RECT  9.520 2.900 9.680 4.140 ;
        RECT  8.840 2.900 9.680 3.100 ;
        RECT  8.980 3.980 9.180 4.400 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.018  LAYER ME1  ;
        ANTENNADIFFAREA 0.978  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.020 2.720 10.300 4.420 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.620 0.900 5.160 1.220 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.100 2.760 1.500 3.160 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 3.680 2.560 3.840 ;
        RECT  2.400 3.420 2.560 3.840 ;
        RECT  0.500 3.920 1.720 4.080 ;
        RECT  1.560 3.680 1.720 4.080 ;
        RECT  0.500 3.640 0.700 4.080 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  8.460 2.260 8.660 3.170 ;
        RECT  7.400 2.260 7.600 3.360 ;
        RECT  0.660 1.730 0.940 3.120 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.500 -0.140 9.700 0.610 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.460 -0.140 7.660 0.560 ;
        RECT  4.460 -0.140 4.660 0.420 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 10.400 4.940 ;
        RECT  9.460 4.300 9.740 4.940 ;
        RECT  8.460 4.240 8.660 4.940 ;
        RECT  7.380 4.240 7.580 4.940 ;
        RECT  5.240 4.240 5.440 4.940 ;
        RECT  3.360 4.380 3.520 4.940 ;
        RECT  0.660 4.480 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.660 2.760 1.860 3.480 ;
        RECT  0.140 3.320 1.860 3.480 ;
        RECT  0.140 3.060 0.340 4.480 ;
        RECT  2.060 0.980 2.800 1.140 ;
        RECT  0.960 0.950 1.160 1.570 ;
        RECT  2.060 0.980 2.220 1.570 ;
        RECT  0.140 1.410 2.220 1.570 ;
        RECT  0.140 0.320 0.340 1.910 ;
        RECT  2.520 3.060 2.880 3.260 ;
        RECT  2.720 3.060 2.880 4.180 ;
        RECT  2.140 4.020 2.880 4.180 ;
        RECT  2.060 0.620 3.120 0.780 ;
        RECT  2.960 1.020 3.560 1.220 ;
        RECT  2.960 0.620 3.120 1.460 ;
        RECT  2.380 1.300 3.120 1.460 ;
        RECT  2.380 1.300 2.540 2.070 ;
        RECT  1.620 1.870 2.540 2.070 ;
        RECT  3.620 0.620 3.980 0.780 ;
        RECT  3.780 0.620 3.980 1.780 ;
        RECT  2.920 1.620 3.980 1.780 ;
        RECT  2.920 1.620 3.120 2.080 ;
        RECT  3.660 3.050 4.280 3.250 ;
        RECT  4.000 3.050 4.280 4.180 ;
        RECT  1.140 0.300 4.300 0.460 ;
        RECT  4.140 0.300 4.300 0.740 ;
        RECT  1.140 0.300 1.340 0.600 ;
        RECT  5.040 0.370 5.200 0.740 ;
        RECT  4.140 0.580 5.200 0.740 ;
        RECT  4.140 0.940 4.300 1.740 ;
        RECT  4.140 1.580 5.300 1.740 ;
        RECT  2.040 2.720 5.660 2.880 ;
        RECT  5.460 2.720 5.660 3.110 ;
        RECT  2.040 2.720 2.240 3.190 ;
        RECT  4.920 3.920 5.920 4.080 ;
        RECT  3.040 4.060 3.840 4.220 ;
        RECT  3.680 4.060 3.840 4.500 ;
        RECT  5.720 3.920 5.920 4.430 ;
        RECT  3.040 4.060 3.200 4.500 ;
        RECT  1.540 4.340 3.200 4.500 ;
        RECT  4.920 3.920 5.080 4.500 ;
        RECT  3.680 4.340 5.080 4.500 ;
        RECT  4.980 3.060 5.180 3.600 ;
        RECT  4.480 3.440 6.620 3.600 ;
        RECT  6.460 3.440 6.620 4.020 ;
        RECT  4.480 3.440 4.760 4.180 ;
        RECT  5.980 2.720 6.940 2.920 ;
        RECT  5.980 2.720 6.180 3.110 ;
        RECT  6.780 2.720 6.940 4.460 ;
        RECT  6.220 4.300 6.940 4.460 ;
        RECT  6.700 1.300 7.680 1.500 ;
        RECT  6.700 0.660 6.980 1.750 ;
        RECT  6.020 0.340 7.300 0.500 ;
        RECT  7.140 0.340 7.300 1.140 ;
        RECT  7.140 0.980 8.240 1.140 ;
        RECT  8.040 0.980 8.240 1.260 ;
        RECT  6.020 0.340 6.180 1.730 ;
        RECT  6.020 1.570 6.500 1.730 ;
        RECT  7.940 0.390 8.140 0.820 ;
        RECT  7.940 0.660 8.780 0.820 ;
        RECT  8.620 0.660 8.780 1.660 ;
        RECT  7.860 1.500 8.780 1.660 ;
        RECT  8.980 0.430 9.180 1.720 ;
        RECT  7.940 3.580 9.360 3.780 ;
        RECT  7.940 2.890 8.140 4.420 ;
        RECT  5.460 0.320 5.820 0.520 ;
        RECT  5.620 0.320 5.820 2.100 ;
        RECT  9.660 0.980 9.860 2.100 ;
        RECT  3.320 1.940 9.860 2.100 ;
        RECT  10.020 0.380 10.220 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.850 3.660 ;
        RECT  2.500 1.140 6.400 3.660 ;
        RECT  0.000 1.160 6.400 3.660 ;
        RECT  7.250 1.140 10.400 3.660 ;
        RECT  0.000 1.180 10.400 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 10.400 4.800 ;
        RECT  0.000 0.000 10.400 1.140 ;
        RECT  1.850 0.000 2.500 1.160 ;
        RECT  6.400 0.000 7.250 1.180 ;
    END
END SDFEZRM4HM

MACRO SDFEZRM2HM
    CLASS CORE ;
    FOREIGN SDFEZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 3.570 3.720 3.900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 0.840 1.900 1.210 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 0.720 1.250 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.345  LAYER ME1  ;
        ANTENNADIFFAREA 0.719  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.980 3.940 9.680 4.120 ;
        RECT  9.520 2.900 9.680 4.120 ;
        RECT  8.930 2.900 9.680 3.260 ;
        RECT  8.980 3.940 9.180 4.500 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.842  LAYER ME1  ;
        ANTENNADIFFAREA 0.719  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.020 3.080 10.300 4.500 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.620 0.900 5.160 1.220 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.100 2.760 1.500 3.160 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 3.680 2.560 3.840 ;
        RECT  2.400 3.420 2.560 3.840 ;
        RECT  0.500 3.920 1.720 4.080 ;
        RECT  1.560 3.680 1.720 4.080 ;
        RECT  0.500 3.640 0.700 4.080 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  8.460 2.260 8.660 3.360 ;
        RECT  7.400 2.260 7.600 3.360 ;
        RECT  0.660 1.730 0.940 3.120 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.500 -0.140 9.700 0.580 ;
        RECT  8.420 -0.140 8.700 0.520 ;
        RECT  7.460 -0.140 7.660 0.560 ;
        RECT  4.460 -0.140 4.660 0.420 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 10.400 4.940 ;
        RECT  9.460 4.280 9.740 4.940 ;
        RECT  8.460 4.220 8.660 4.940 ;
        RECT  7.380 4.240 7.580 4.940 ;
        RECT  5.240 4.240 5.440 4.940 ;
        RECT  3.360 4.380 3.520 4.940 ;
        RECT  0.660 4.480 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.660 2.760 1.860 3.480 ;
        RECT  0.140 3.320 1.860 3.480 ;
        RECT  0.140 3.060 0.340 4.480 ;
        RECT  2.060 0.980 2.800 1.140 ;
        RECT  0.960 0.950 1.160 1.570 ;
        RECT  2.060 0.980 2.220 1.570 ;
        RECT  0.140 1.410 2.220 1.570 ;
        RECT  0.140 0.320 0.340 1.910 ;
        RECT  2.520 3.060 2.880 3.260 ;
        RECT  2.720 3.060 2.880 4.180 ;
        RECT  2.140 4.020 2.880 4.180 ;
        RECT  2.060 0.620 3.120 0.780 ;
        RECT  2.960 1.020 3.560 1.220 ;
        RECT  2.960 0.620 3.120 1.460 ;
        RECT  2.380 1.300 3.120 1.460 ;
        RECT  2.380 1.300 2.540 2.070 ;
        RECT  1.620 1.870 2.540 2.070 ;
        RECT  3.620 0.620 3.980 0.780 ;
        RECT  3.780 0.620 3.980 1.780 ;
        RECT  2.920 1.620 3.980 1.780 ;
        RECT  2.920 1.620 3.120 2.080 ;
        RECT  3.660 3.050 4.280 3.250 ;
        RECT  4.000 3.050 4.280 4.180 ;
        RECT  1.140 0.300 4.300 0.460 ;
        RECT  4.140 0.300 4.300 0.740 ;
        RECT  1.140 0.300 1.340 0.600 ;
        RECT  5.040 0.370 5.200 0.740 ;
        RECT  4.140 0.580 5.200 0.740 ;
        RECT  4.140 0.940 4.300 1.740 ;
        RECT  4.140 1.580 5.300 1.740 ;
        RECT  2.040 2.720 5.660 2.880 ;
        RECT  5.460 2.720 5.660 3.110 ;
        RECT  2.040 2.720 2.240 3.190 ;
        RECT  4.920 3.920 5.920 4.080 ;
        RECT  3.040 4.060 3.840 4.220 ;
        RECT  3.680 4.060 3.840 4.500 ;
        RECT  5.720 3.920 5.920 4.430 ;
        RECT  3.040 4.060 3.200 4.500 ;
        RECT  1.540 4.340 3.200 4.500 ;
        RECT  4.920 3.920 5.080 4.500 ;
        RECT  3.680 4.340 5.080 4.500 ;
        RECT  4.980 3.060 5.180 3.600 ;
        RECT  4.480 3.440 6.620 3.600 ;
        RECT  6.460 3.440 6.620 4.020 ;
        RECT  4.480 3.440 4.760 4.180 ;
        RECT  5.980 2.720 6.940 2.920 ;
        RECT  5.980 2.720 6.180 3.110 ;
        RECT  6.780 2.720 6.940 4.460 ;
        RECT  6.220 4.300 6.940 4.460 ;
        RECT  6.700 1.320 7.720 1.480 ;
        RECT  6.700 0.660 6.980 1.750 ;
        RECT  6.020 0.340 7.300 0.500 ;
        RECT  7.140 0.340 7.300 1.160 ;
        RECT  7.140 1.000 8.240 1.160 ;
        RECT  8.040 1.000 8.240 1.280 ;
        RECT  6.020 0.340 6.180 1.730 ;
        RECT  6.020 1.570 6.500 1.730 ;
        RECT  7.940 0.390 8.140 0.840 ;
        RECT  7.940 0.680 8.780 0.840 ;
        RECT  8.620 0.680 8.780 1.780 ;
        RECT  7.900 1.580 8.780 1.780 ;
        RECT  8.980 0.300 9.180 1.720 ;
        RECT  7.940 3.580 9.360 3.780 ;
        RECT  7.940 3.000 8.140 4.440 ;
        RECT  5.460 0.320 5.820 0.520 ;
        RECT  5.620 0.320 5.820 2.100 ;
        RECT  9.660 0.980 9.860 2.100 ;
        RECT  3.320 1.940 9.860 2.100 ;
        RECT  10.020 0.300 10.220 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.850 3.660 ;
        RECT  2.500 1.140 6.400 3.660 ;
        RECT  0.000 1.160 6.400 3.660 ;
        RECT  7.250 1.140 10.400 3.660 ;
        RECT  0.000 1.180 10.400 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 10.400 4.800 ;
        RECT  0.000 0.000 10.400 1.140 ;
        RECT  1.850 0.000 2.500 1.160 ;
        RECT  6.400 0.000 7.250 1.180 ;
    END
END SDFEZRM2HM

MACRO SDFEZRM1HM
    CLASS CORE ;
    FOREIGN SDFEZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        ANTENNAGATEAREA 0.161  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.694  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.030 0.940 7.230 1.140 ;
        LAYER ME1 ;
        RECT  6.940 0.920 8.790 1.080 ;
        RECT  6.940 0.920 7.370 1.140 ;
        LAYER ME2 ;
        RECT  6.900 0.750 7.230 1.250 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.047  LAYER ME1  ;
        ANTENNAGATEAREA 0.047  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.556  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.340 6.300 1.540 ;
        LAYER ME1 ;
        RECT  5.830 1.340 6.400 1.540 ;
        LAYER ME2 ;
        RECT  6.100 1.100 6.300 1.690 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.200 1.050 9.500 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.610 1.190 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.430 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.319  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.010 0.840 17.500 1.160 ;
        RECT  17.010 0.350 17.230 1.760 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  18.230 1.650 18.700 1.850 ;
        RECT  18.500 0.370 18.700 1.850 ;
        RECT  18.230 0.370 18.700 0.570 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 0.840 3.520 1.310 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.800 2.540 ;
        RECT  17.710 1.640 17.910 2.540 ;
        RECT  15.910 2.020 16.110 2.540 ;
        RECT  12.620 1.860 12.900 2.540 ;
        RECT  8.860 2.080 9.140 2.540 ;
        RECT  5.870 2.020 6.070 2.540 ;
        RECT  4.140 1.520 4.340 2.540 ;
        RECT  3.060 1.860 3.340 2.540 ;
        RECT  2.420 1.860 2.700 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.800 0.140 ;
        RECT  17.710 -0.140 17.910 0.610 ;
        RECT  15.870 -0.140 16.070 0.560 ;
        RECT  12.620 -0.140 12.900 0.320 ;
        RECT  8.410 -0.140 8.610 0.380 ;
        RECT  6.090 -0.140 6.370 0.540 ;
        RECT  3.780 -0.140 3.980 0.560 ;
        RECT  0.100 -0.140 0.380 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.370 1.000 0.570 ;
        RECT  1.770 1.040 2.520 1.240 ;
        RECT  0.800 0.370 1.000 1.700 ;
        RECT  0.140 1.510 1.000 1.700 ;
        RECT  1.770 1.040 1.930 1.700 ;
        RECT  0.140 1.540 1.930 1.700 ;
        RECT  0.140 1.510 0.340 1.870 ;
        RECT  1.160 0.300 3.380 0.460 ;
        RECT  1.160 0.300 1.360 0.600 ;
        RECT  3.180 0.300 3.380 0.620 ;
        RECT  2.220 0.620 2.840 0.780 ;
        RECT  3.780 0.960 4.360 1.170 ;
        RECT  2.680 0.620 2.840 1.700 ;
        RECT  3.780 0.960 3.940 1.700 ;
        RECT  2.090 1.540 3.940 1.700 ;
        RECT  2.090 1.540 2.250 2.020 ;
        RECT  1.540 1.860 2.250 2.020 ;
        RECT  4.670 0.300 5.930 0.460 ;
        RECT  6.530 0.300 7.390 0.500 ;
        RECT  4.260 0.400 4.870 0.600 ;
        RECT  5.770 0.300 5.930 0.860 ;
        RECT  6.530 0.300 6.690 0.860 ;
        RECT  5.770 0.700 6.690 0.860 ;
        RECT  4.670 0.300 4.870 1.700 ;
        RECT  5.320 0.620 5.600 1.180 ;
        RECT  5.190 1.020 6.750 1.180 ;
        RECT  7.780 1.240 8.060 1.460 ;
        RECT  6.590 1.300 8.060 1.460 ;
        RECT  6.590 1.020 6.750 1.630 ;
        RECT  5.190 1.020 5.390 1.780 ;
        RECT  8.220 1.400 8.690 1.600 ;
        RECT  8.220 1.400 8.380 1.780 ;
        RECT  6.910 1.620 8.380 1.780 ;
        RECT  9.090 0.620 9.880 0.780 ;
        RECT  9.680 0.830 10.230 1.030 ;
        RECT  9.680 0.620 9.880 1.780 ;
        RECT  10.520 0.620 10.880 0.840 ;
        RECT  10.680 1.080 11.000 1.360 ;
        RECT  10.680 0.620 10.880 1.780 ;
        RECT  8.770 0.300 11.240 0.460 ;
        RECT  7.550 0.350 7.710 0.710 ;
        RECT  11.040 0.300 11.240 0.610 ;
        RECT  8.770 0.300 8.930 0.710 ;
        RECT  7.550 0.550 8.930 0.710 ;
        RECT  11.080 1.500 11.480 1.780 ;
        RECT  11.580 0.380 11.740 1.200 ;
        RECT  11.740 1.220 13.150 1.380 ;
        RECT  11.740 1.040 11.940 1.780 ;
        RECT  13.380 0.620 13.660 0.960 ;
        RECT  12.360 0.800 13.660 0.960 ;
        RECT  13.460 0.620 13.660 1.740 ;
        RECT  13.460 1.540 13.870 1.740 ;
        RECT  13.060 0.300 13.980 0.460 ;
        RECT  13.060 0.300 13.220 0.640 ;
        RECT  11.940 0.480 13.220 0.640 ;
        RECT  11.940 0.480 12.140 0.860 ;
        RECT  13.820 0.300 13.980 1.150 ;
        RECT  14.150 0.300 15.670 0.460 ;
        RECT  15.510 0.300 15.670 1.160 ;
        RECT  15.510 1.000 16.290 1.160 ;
        RECT  14.150 0.300 14.350 1.780 ;
        RECT  16.450 1.020 16.790 1.300 ;
        RECT  16.450 0.430 16.650 1.480 ;
        RECT  15.370 1.320 16.750 1.480 ;
        RECT  16.590 1.020 16.750 1.780 ;
        RECT  14.770 0.620 15.350 0.780 ;
        RECT  17.930 0.960 18.130 1.480 ;
        RECT  17.390 1.320 18.130 1.480 ;
        RECT  12.100 1.540 13.220 1.700 ;
        RECT  5.550 1.700 6.390 1.860 ;
        RECT  14.770 1.700 16.430 1.860 ;
        RECT  8.540 1.760 9.460 1.920 ;
        RECT  6.230 1.700 6.390 2.100 ;
        RECT  9.300 1.760 9.460 2.100 ;
        RECT  13.060 1.540 13.220 2.100 ;
        RECT  16.270 1.700 16.430 2.100 ;
        RECT  5.550 1.700 5.710 2.100 ;
        RECT  4.780 1.940 5.710 2.100 ;
        RECT  8.540 1.760 8.700 2.100 ;
        RECT  6.230 1.940 8.700 2.100 ;
        RECT  12.100 1.540 12.260 2.100 ;
        RECT  9.300 1.940 12.260 2.100 ;
        RECT  14.770 0.620 14.930 2.100 ;
        RECT  13.060 1.940 14.930 2.100 ;
        RECT  17.390 1.320 17.550 2.100 ;
        RECT  16.270 1.940 17.550 2.100 ;
        LAYER VI1 ;
        RECT  8.390 1.400 8.590 1.600 ;
        RECT  11.180 1.580 11.380 1.780 ;
        LAYER ME2 ;
        RECT  8.390 1.300 8.590 1.960 ;
        RECT  11.180 1.480 11.380 1.960 ;
        RECT  8.390 1.760 11.380 1.960 ;
        LAYER VTPH ;
        RECT  0.420 1.030 2.020 2.400 ;
        RECT  3.760 1.010 5.070 2.400 ;
        RECT  11.060 1.000 12.100 2.400 ;
        RECT  0.000 1.140 18.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.800 1.000 ;
        RECT  0.000 0.000 11.060 1.010 ;
        RECT  0.000 0.000 3.760 1.030 ;
        RECT  0.000 0.000 0.420 1.140 ;
        RECT  2.020 0.000 3.760 1.140 ;
        RECT  5.070 0.000 11.060 1.140 ;
        RECT  12.100 0.000 18.800 1.140 ;
    END
END SDFEZRM1HM

MACRO SDFERM8HM
    CLASS CORE ;
    FOREIGN SDFERM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        ANTENNAGATEAREA 0.199  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.141  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.360 1.110 7.560 1.310 ;
        LAYER ME2 ;
        RECT  7.300 0.840 7.560 1.560 ;
        LAYER ME1 ;
        RECT  7.360 0.900 7.620 1.460 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.108  LAYER ME1  ;
        ANTENNAGATEAREA 0.108  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.659  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.850 1.070 5.050 1.270 ;
        LAYER ME2 ;
        RECT  4.810 0.840 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.720 0.950 5.080 1.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.133  LAYER ME1  ;
        ANTENNAGATEAREA 0.133  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.162  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.970 1.050 8.170 1.250 ;
        LAYER ME2 ;
        RECT  7.970 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  7.800 0.900 8.170 1.340 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.968  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 3.040 2.440 3.300 ;
        RECT  2.240 3.960 2.400 4.390 ;
        RECT  1.200 3.960 2.400 4.120 ;
        RECT  1.200 3.040 1.360 4.460 ;
        RECT  0.900 3.040 1.360 3.750 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.874  LAYER ME1  ;
        ANTENNADIFFAREA 1.394  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.520 1.360 1.680 ;
        RECT  0.100 0.690 1.360 0.860 ;
        RECT  1.200 0.330 1.360 0.860 ;
        RECT  0.100 0.690 0.330 1.680 ;
        RECT  0.100 0.360 0.320 2.070 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.386  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 3.550 4.300 3.750 ;
        LAYER ME2 ;
        RECT  4.100 3.240 4.300 3.960 ;
        LAYER ME1 ;
        RECT  4.040 3.540 4.740 3.750 ;
        RECT  4.040 3.340 4.360 3.750 ;
        RECT  2.930 3.340 4.360 3.500 ;
        RECT  2.930 3.340 3.090 3.790 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.425  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.780 3.900 0.980 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  3.540 0.710 4.080 1.040 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.163  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.260 1.100 4.460 1.300 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.460 1.560 ;
        LAYER ME1 ;
        RECT  2.970 1.200 4.560 1.360 ;
        RECT  4.260 1.030 4.560 1.360 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.020 1.570 10.310 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  7.690 -0.140 7.850 0.420 ;
        RECT  1.700 -0.140 1.980 0.380 ;
        RECT  0.600 -0.140 0.920 0.500 ;
        RECT  0.000 4.660 11.200 4.940 ;
        RECT  7.930 4.260 8.210 4.940 ;
        RECT  4.600 4.260 4.880 4.940 ;
        RECT  2.700 4.270 2.980 4.940 ;
        RECT  1.660 4.280 1.940 4.940 ;
        RECT  0.680 4.080 0.840 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 2.860 0.320 4.380 ;
        RECT  0.490 1.020 1.580 1.240 ;
        RECT  2.480 0.740 3.260 0.900 ;
        RECT  1.830 1.080 2.640 1.240 ;
        RECT  2.480 0.740 2.640 1.780 ;
        RECT  2.480 1.550 4.560 1.780 ;
        RECT  2.600 3.020 5.120 3.180 ;
        RECT  1.540 3.570 2.770 3.730 ;
        RECT  4.960 3.020 5.120 3.740 ;
        RECT  2.600 3.020 2.770 4.110 ;
        RECT  2.600 3.950 3.300 4.110 ;
        RECT  3.140 3.950 3.300 4.450 ;
        RECT  3.140 4.290 3.960 4.450 ;
        RECT  0.500 2.700 5.590 2.860 ;
        RECT  5.280 2.700 5.590 2.920 ;
        RECT  5.280 2.700 5.520 3.400 ;
        RECT  0.500 2.700 0.660 3.880 ;
        RECT  5.360 2.700 5.520 4.180 ;
        RECT  5.360 3.910 5.640 4.180 ;
        RECT  2.160 0.300 5.870 0.460 ;
        RECT  5.570 0.300 5.870 0.570 ;
        RECT  2.160 0.300 2.320 0.800 ;
        RECT  1.960 0.640 2.320 0.800 ;
        RECT  2.060 1.780 2.300 2.100 ;
        RECT  5.630 1.890 5.970 2.100 ;
        RECT  2.060 1.940 5.970 2.100 ;
        RECT  6.100 3.020 6.600 3.260 ;
        RECT  3.460 3.660 3.740 4.100 ;
        RECT  3.460 3.940 5.200 4.100 ;
        RECT  5.040 3.940 5.200 4.500 ;
        RECT  5.920 3.980 6.260 4.500 ;
        RECT  6.100 3.020 6.260 4.500 ;
        RECT  5.040 4.340 6.260 4.500 ;
        RECT  5.480 1.070 7.200 1.230 ;
        RECT  5.480 1.070 5.770 1.390 ;
        RECT  7.000 0.620 7.200 1.780 ;
        RECT  7.000 1.620 7.400 1.780 ;
        RECT  7.250 3.020 8.770 3.220 ;
        RECT  8.490 3.020 8.770 3.460 ;
        RECT  7.250 3.020 7.410 4.180 ;
        RECT  6.820 3.850 7.410 4.180 ;
        RECT  4.720 1.550 6.290 1.710 ;
        RECT  4.720 1.550 5.080 1.780 ;
        RECT  6.130 1.550 6.290 2.100 ;
        RECT  6.130 1.940 8.890 2.100 ;
        RECT  7.610 3.940 9.420 4.100 ;
        RECT  6.420 3.420 6.580 4.500 ;
        RECT  7.610 3.940 7.770 4.500 ;
        RECT  6.420 4.340 7.770 4.500 ;
        RECT  8.330 0.640 8.610 1.180 ;
        RECT  8.330 1.020 9.510 1.180 ;
        RECT  8.330 0.640 8.490 1.760 ;
        RECT  8.070 1.500 8.490 1.760 ;
        RECT  7.590 3.500 7.890 3.780 ;
        RECT  7.590 3.620 10.230 3.780 ;
        RECT  9.950 3.340 10.230 4.420 ;
        RECT  9.780 3.620 10.230 4.420 ;
        RECT  6.520 0.300 7.530 0.460 ;
        RECT  8.010 0.300 10.200 0.460 ;
        RECT  7.370 0.300 7.530 0.740 ;
        RECT  10.040 0.300 10.200 0.740 ;
        RECT  8.010 0.300 8.170 0.740 ;
        RECT  7.370 0.580 8.170 0.740 ;
        RECT  10.040 0.580 10.480 0.740 ;
        RECT  4.510 0.620 5.410 0.780 ;
        RECT  6.520 0.300 6.760 0.910 ;
        RECT  5.250 0.750 6.760 0.910 ;
        RECT  5.780 2.700 10.540 2.860 ;
        RECT  6.880 2.700 7.080 3.670 ;
        RECT  5.780 2.700 5.940 3.740 ;
        RECT  5.680 3.340 5.940 3.740 ;
        RECT  8.930 3.020 10.770 3.180 ;
        RECT  8.930 3.020 9.130 3.310 ;
        RECT  10.570 3.020 10.770 3.380 ;
        RECT  9.290 0.620 9.860 0.780 ;
        RECT  9.700 1.250 10.830 1.410 ;
        RECT  9.700 0.620 9.860 1.680 ;
        RECT  8.670 1.460 9.860 1.680 ;
        RECT  10.520 1.250 10.830 1.690 ;
        RECT  10.760 3.570 10.920 4.380 ;
        RECT  10.520 4.220 10.920 4.380 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.880 3.660 ;
        RECT  0.000 1.160 2.520 3.660 ;
        RECT  4.410 1.210 5.620 3.600 ;
        RECT  7.450 1.160 11.200 3.540 ;
        RECT  0.000 1.260 11.200 3.540 ;
        RECT  0.000 1.260 5.780 3.600 ;
        RECT  0.000 1.260 4.470 3.660 ;
        RECT  9.870 1.140 11.200 3.660 ;
        RECT  8.630 1.160 10.660 3.860 ;
        LAYER VTNH ;
        RECT  4.470 3.600 8.630 4.800 ;
        RECT  5.780 3.540 8.630 4.800 ;
        RECT  0.000 3.660 8.630 4.800 ;
        RECT  10.660 3.660 11.200 4.800 ;
        RECT  0.000 3.860 11.200 4.800 ;
        RECT  0.000 0.000 11.200 1.140 ;
        RECT  1.880 0.000 9.870 1.160 ;
        RECT  2.520 0.000 7.450 1.210 ;
        RECT  2.520 0.000 4.410 1.260 ;
        RECT  5.620 0.000 7.450 1.260 ;
    END
END SDFERM8HM

MACRO SDFERM4HM
    CLASS CORE ;
    FOREIGN SDFERM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.108  LAYER ME1  ;
        ANTENNAGATEAREA 0.108  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.659  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.070 3.900 1.270 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.690 0.950 4.050 1.350 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        ANTENNAGATEAREA 0.199  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.141  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.330 1.110 6.530 1.310 ;
        LAYER ME2 ;
        RECT  6.100 0.840 6.530 1.560 ;
        LAYER ME1 ;
        RECT  6.330 0.900 6.590 1.460 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.770 0.900 7.210 1.340 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.498  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 3.040 1.460 3.300 ;
        RECT  1.260 3.960 1.420 4.390 ;
        RECT  0.900 3.960 1.420 4.120 ;
        RECT  0.900 3.040 1.100 4.120 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.924  LAYER ME1  ;
        ANTENNADIFFAREA 0.843  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.750 0.320 2.070 ;
        RECT  0.100 0.360 0.320 0.730 ;
        RECT  0.100 0.360 0.300 2.070 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.985  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.250 3.550 3.450 3.750 ;
        LAYER ME2 ;
        RECT  3.250 3.240 3.500 3.960 ;
        LAYER ME1 ;
        RECT  3.020 3.340 3.540 3.750 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.183  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 0.780 2.700 0.980 ;
        LAYER ME2 ;
        RECT  2.500 0.440 2.700 1.160 ;
        LAYER ME1 ;
        RECT  2.440 0.710 3.050 1.040 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.163  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.100 3.500 1.300 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  1.940 1.200 3.530 1.360 ;
        RECT  3.230 1.030 3.530 1.360 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  8.820 1.570 9.110 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  6.660 -0.140 6.820 0.420 ;
        RECT  0.670 -0.140 0.950 0.380 ;
        RECT  0.000 4.660 10.000 4.940 ;
        RECT  6.730 4.260 7.010 4.940 ;
        RECT  3.340 4.260 3.620 4.940 ;
        RECT  1.720 4.270 2.000 4.940 ;
        RECT  0.630 4.280 0.910 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 2.790 0.320 4.380 ;
        RECT  1.490 0.740 2.270 0.900 ;
        RECT  0.840 1.080 1.650 1.240 ;
        RECT  1.490 0.740 1.650 1.780 ;
        RECT  1.450 1.080 1.650 1.780 ;
        RECT  1.450 1.550 3.530 1.780 ;
        RECT  2.230 3.020 3.860 3.180 ;
        RECT  3.700 3.020 3.860 3.740 ;
        RECT  2.230 3.020 2.400 3.790 ;
        RECT  1.350 3.510 2.400 3.790 ;
        RECT  2.240 3.020 2.400 4.450 ;
        RECT  2.240 4.290 2.700 4.450 ;
        RECT  0.510 2.700 4.330 2.860 ;
        RECT  4.020 2.700 4.330 2.920 ;
        RECT  4.020 2.700 4.260 3.400 ;
        RECT  0.510 2.700 0.670 3.880 ;
        RECT  4.100 2.700 4.260 4.180 ;
        RECT  4.100 3.910 4.380 4.180 ;
        RECT  1.170 0.300 4.840 0.460 ;
        RECT  4.540 0.300 4.840 0.570 ;
        RECT  1.170 0.300 1.330 0.860 ;
        RECT  0.990 0.580 1.330 0.860 ;
        RECT  1.030 1.780 1.270 2.100 ;
        RECT  4.600 1.890 4.940 2.100 ;
        RECT  1.030 1.940 4.940 2.100 ;
        RECT  4.840 3.020 5.340 3.260 ;
        RECT  2.560 3.450 2.760 4.100 ;
        RECT  2.560 3.940 3.940 4.100 ;
        RECT  3.780 3.940 3.940 4.500 ;
        RECT  4.660 3.980 5.000 4.500 ;
        RECT  4.840 3.020 5.000 4.500 ;
        RECT  3.780 4.340 5.000 4.500 ;
        RECT  4.450 1.070 6.170 1.230 ;
        RECT  4.450 1.070 4.740 1.390 ;
        RECT  5.970 0.620 6.170 1.780 ;
        RECT  5.970 1.620 6.370 1.780 ;
        RECT  6.050 3.020 7.570 3.220 ;
        RECT  7.290 3.020 7.570 3.460 ;
        RECT  6.050 3.020 6.210 4.180 ;
        RECT  5.830 3.880 6.210 4.180 ;
        RECT  3.690 1.550 5.260 1.710 ;
        RECT  3.690 1.550 4.050 1.780 ;
        RECT  5.100 1.550 5.260 2.100 ;
        RECT  5.100 1.940 8.080 2.100 ;
        RECT  6.410 3.940 8.220 4.100 ;
        RECT  5.160 3.420 5.320 4.500 ;
        RECT  6.410 3.940 6.570 4.500 ;
        RECT  5.160 4.340 6.570 4.500 ;
        RECT  7.370 0.640 7.650 1.240 ;
        RECT  7.370 0.960 8.250 1.240 ;
        RECT  7.370 0.640 7.530 1.760 ;
        RECT  7.110 1.500 7.530 1.760 ;
        RECT  6.390 3.500 6.690 3.780 ;
        RECT  6.390 3.620 9.030 3.780 ;
        RECT  8.750 3.340 9.030 4.420 ;
        RECT  8.580 3.620 9.030 4.420 ;
        RECT  4.520 2.700 9.340 2.860 ;
        RECT  5.620 2.700 5.820 3.690 ;
        RECT  4.520 2.700 4.680 3.740 ;
        RECT  4.420 3.340 4.680 3.740 ;
        RECT  7.730 3.020 9.570 3.180 ;
        RECT  7.730 3.020 7.930 3.310 ;
        RECT  9.370 3.020 9.570 3.380 ;
        RECT  5.490 0.300 6.500 0.460 ;
        RECT  6.980 0.300 9.290 0.460 ;
        RECT  6.340 0.300 6.500 0.740 ;
        RECT  9.130 0.300 9.290 0.740 ;
        RECT  6.980 0.300 7.140 0.740 ;
        RECT  6.340 0.580 7.140 0.740 ;
        RECT  9.130 0.580 9.570 0.740 ;
        RECT  3.480 0.620 4.380 0.780 ;
        RECT  5.490 0.300 5.730 0.910 ;
        RECT  4.220 0.750 5.730 0.910 ;
        RECT  8.310 0.620 8.650 0.780 ;
        RECT  8.410 0.620 8.650 1.410 ;
        RECT  8.410 1.250 9.630 1.410 ;
        RECT  9.320 1.250 9.630 1.690 ;
        RECT  8.410 0.620 8.590 1.710 ;
        RECT  7.860 1.490 8.590 1.710 ;
        RECT  9.560 3.570 9.720 4.380 ;
        RECT  9.320 4.220 9.720 4.380 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.890 3.660 ;
        RECT  0.000 1.160 1.530 3.660 ;
        RECT  3.380 1.210 4.590 3.540 ;
        RECT  6.420 1.160 10.000 3.540 ;
        RECT  0.000 1.260 10.000 3.540 ;
        RECT  0.000 1.260 4.520 3.600 ;
        RECT  0.000 1.260 3.210 3.660 ;
        RECT  8.780 1.140 10.000 3.660 ;
        RECT  7.430 1.160 9.460 3.860 ;
        LAYER VTNH ;
        RECT  3.210 3.600 7.430 4.800 ;
        RECT  4.520 3.540 7.430 4.800 ;
        RECT  0.000 3.660 7.430 4.800 ;
        RECT  9.460 3.660 10.000 4.800 ;
        RECT  0.000 3.860 10.000 4.800 ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  0.890 0.000 8.780 1.160 ;
        RECT  1.530 0.000 6.420 1.210 ;
        RECT  1.530 0.000 3.380 1.260 ;
        RECT  4.590 0.000 6.420 1.260 ;
    END
END SDFERM4HM

MACRO SDFERM2HM
    CLASS CORE ;
    FOREIGN SDFERM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        ANTENNAGATEAREA 0.199  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.141  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.930 1.110 6.130 1.310 ;
        LAYER ME2 ;
        RECT  5.700 0.840 6.130 1.560 ;
        LAYER ME1 ;
        RECT  5.930 0.900 6.190 1.460 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.108  LAYER ME1  ;
        ANTENNAGATEAREA 0.108  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.659  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.070 3.500 1.270 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.290 0.950 3.650 1.350 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.536  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.850 3.550 3.050 3.750 ;
        LAYER ME2 ;
        RECT  2.850 3.240 3.100 3.960 ;
        LAYER ME1 ;
        RECT  2.760 3.340 3.140 3.750 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.370 0.900 6.810 1.340 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.433  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 3.040 1.670 4.390 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 2.720 0.340 4.380 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.183  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 0.780 2.300 0.980 ;
        LAYER ME2 ;
        RECT  2.100 0.440 2.300 1.160 ;
        LAYER ME1 ;
        RECT  2.040 0.710 2.650 1.040 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.172  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.100 3.100 1.300 ;
        LAYER ME2 ;
        RECT  2.900 0.840 3.100 1.560 ;
        LAYER ME1 ;
        RECT  1.540 1.200 3.130 1.360 ;
        RECT  2.830 1.030 3.130 1.360 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.420 1.570 8.710 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  6.260 -0.140 6.420 0.420 ;
        RECT  0.100 -0.140 0.380 0.380 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  6.330 4.260 6.610 4.940 ;
        RECT  2.940 4.260 3.220 4.940 ;
        RECT  0.800 4.270 1.080 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.090 0.740 1.770 0.900 ;
        RECT  0.220 1.060 1.250 1.260 ;
        RECT  1.090 0.740 1.250 1.780 ;
        RECT  1.050 1.060 1.250 1.780 ;
        RECT  1.050 1.550 3.130 1.780 ;
        RECT  1.990 3.020 3.460 3.180 ;
        RECT  3.300 3.020 3.460 3.740 ;
        RECT  1.990 3.020 2.160 3.790 ;
        RECT  1.860 3.510 2.160 3.790 ;
        RECT  2.000 3.020 2.160 4.500 ;
        RECT  2.000 4.260 2.300 4.500 ;
        RECT  0.560 2.700 3.930 2.860 ;
        RECT  3.620 2.700 3.930 2.920 ;
        RECT  3.620 2.700 3.860 3.400 ;
        RECT  0.560 2.700 0.780 3.880 ;
        RECT  3.700 2.700 3.860 4.180 ;
        RECT  3.700 3.910 3.980 4.180 ;
        RECT  0.770 0.300 4.440 0.460 ;
        RECT  4.140 0.300 4.440 0.570 ;
        RECT  0.770 0.300 0.930 0.860 ;
        RECT  0.420 0.580 0.930 0.860 ;
        RECT  0.420 1.690 0.660 2.100 ;
        RECT  4.200 1.890 4.540 2.100 ;
        RECT  0.420 1.940 4.540 2.100 ;
        RECT  4.440 3.020 4.940 3.260 ;
        RECT  2.320 3.450 2.520 4.100 ;
        RECT  2.320 3.940 3.540 4.100 ;
        RECT  3.380 3.940 3.540 4.500 ;
        RECT  4.260 3.980 4.600 4.500 ;
        RECT  4.440 3.020 4.600 4.500 ;
        RECT  3.380 4.340 4.600 4.500 ;
        RECT  4.050 1.070 5.770 1.230 ;
        RECT  4.050 1.070 4.340 1.390 ;
        RECT  5.570 0.620 5.770 1.780 ;
        RECT  5.570 1.620 5.970 1.780 ;
        RECT  5.650 3.020 7.170 3.220 ;
        RECT  6.890 3.020 7.170 3.460 ;
        RECT  5.650 3.020 5.810 4.180 ;
        RECT  5.430 3.880 5.810 4.180 ;
        RECT  3.290 1.550 4.860 1.710 ;
        RECT  3.290 1.550 3.650 1.780 ;
        RECT  4.700 1.550 4.860 2.100 ;
        RECT  4.700 1.940 7.680 2.100 ;
        RECT  6.010 3.940 7.820 4.100 ;
        RECT  4.760 3.420 4.920 4.500 ;
        RECT  6.010 3.940 6.170 4.500 ;
        RECT  4.760 4.340 6.170 4.500 ;
        RECT  6.970 0.640 7.250 1.240 ;
        RECT  6.970 0.960 7.850 1.240 ;
        RECT  6.970 0.640 7.130 1.760 ;
        RECT  6.710 1.500 7.130 1.760 ;
        RECT  5.990 3.500 6.290 3.780 ;
        RECT  5.990 3.620 8.630 3.780 ;
        RECT  8.350 3.340 8.630 4.420 ;
        RECT  8.180 3.620 8.630 4.420 ;
        RECT  4.120 2.700 8.940 2.860 ;
        RECT  5.220 2.700 5.420 3.690 ;
        RECT  4.120 2.700 4.280 3.740 ;
        RECT  4.020 3.340 4.280 3.740 ;
        RECT  7.330 3.020 9.170 3.180 ;
        RECT  7.330 3.020 7.530 3.310 ;
        RECT  8.970 3.020 9.170 3.380 ;
        RECT  5.090 0.300 6.100 0.460 ;
        RECT  6.580 0.300 8.890 0.460 ;
        RECT  5.940 0.300 6.100 0.740 ;
        RECT  8.730 0.300 8.890 0.740 ;
        RECT  6.580 0.300 6.740 0.740 ;
        RECT  5.940 0.580 6.740 0.740 ;
        RECT  8.730 0.580 9.170 0.740 ;
        RECT  3.080 0.620 3.980 0.780 ;
        RECT  5.090 0.300 5.330 0.910 ;
        RECT  3.820 0.750 5.330 0.910 ;
        RECT  7.910 0.620 8.250 0.780 ;
        RECT  8.010 0.620 8.250 1.410 ;
        RECT  8.010 1.250 9.230 1.410 ;
        RECT  8.920 1.250 9.230 1.690 ;
        RECT  8.010 0.620 8.190 1.710 ;
        RECT  7.460 1.490 8.190 1.710 ;
        RECT  9.160 3.570 9.320 4.380 ;
        RECT  8.920 4.220 9.320 4.380 ;
        LAYER VTPH ;
        RECT  0.000 1.160 1.130 3.660 ;
        RECT  2.980 1.210 4.190 3.540 ;
        RECT  6.020 1.160 9.600 3.540 ;
        RECT  0.000 1.260 9.600 3.540 ;
        RECT  0.000 1.260 4.120 3.600 ;
        RECT  0.000 1.260 2.810 3.660 ;
        RECT  8.380 1.140 9.600 3.660 ;
        RECT  7.030 1.160 9.060 3.860 ;
        LAYER VTNH ;
        RECT  2.810 3.600 7.030 4.800 ;
        RECT  4.120 3.540 7.030 4.800 ;
        RECT  0.000 3.660 7.030 4.800 ;
        RECT  9.060 3.660 9.600 4.800 ;
        RECT  0.000 3.860 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  0.000 0.000 8.380 1.160 ;
        RECT  1.130 0.000 6.020 1.210 ;
        RECT  1.130 0.000 2.980 1.260 ;
        RECT  4.190 0.000 6.020 1.260 ;
    END
END SDFERM2HM

MACRO SDFERM1HM
    CLASS CORE ;
    FOREIGN SDFERM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        ANTENNAGATEAREA 0.199  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.141  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.930 1.110 6.130 1.310 ;
        LAYER ME2 ;
        RECT  5.700 0.840 6.130 1.560 ;
        LAYER ME1 ;
        RECT  5.930 0.900 6.190 1.460 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.742  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.070 3.500 1.270 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.290 0.950 3.650 1.350 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.458  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.850 3.550 3.050 3.750 ;
        LAYER ME2 ;
        RECT  2.850 3.240 3.100 3.960 ;
        LAYER ME1 ;
        RECT  2.760 3.340 3.140 3.750 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.370 0.900 6.810 1.340 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.304  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 3.040 1.630 4.460 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.340  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 3.080 0.340 4.450 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.183  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 0.780 2.300 0.980 ;
        LAYER ME2 ;
        RECT  2.100 0.440 2.300 1.160 ;
        LAYER ME1 ;
        RECT  2.040 0.710 2.650 1.040 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.172  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.100 3.100 1.300 ;
        LAYER ME2 ;
        RECT  2.900 0.840 3.100 1.560 ;
        LAYER ME1 ;
        RECT  1.540 1.200 3.130 1.360 ;
        RECT  2.830 1.030 3.130 1.360 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.420 1.570 8.710 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  6.260 -0.140 6.420 0.420 ;
        RECT  0.100 -0.140 0.380 0.380 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  6.330 4.260 6.610 4.940 ;
        RECT  2.940 4.260 3.220 4.940 ;
        RECT  0.800 4.270 1.080 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.090 0.740 1.770 0.900 ;
        RECT  0.220 1.060 1.250 1.260 ;
        RECT  1.090 0.740 1.250 1.780 ;
        RECT  1.050 1.060 1.250 1.780 ;
        RECT  1.050 1.550 3.130 1.780 ;
        RECT  1.870 3.020 3.460 3.180 ;
        RECT  3.300 3.020 3.460 3.740 ;
        RECT  1.870 3.020 2.120 3.790 ;
        RECT  1.820 3.510 2.120 3.790 ;
        RECT  1.880 3.020 2.120 4.500 ;
        RECT  1.880 4.260 2.160 4.500 ;
        RECT  0.560 2.700 3.930 2.860 ;
        RECT  3.620 2.700 3.930 2.920 ;
        RECT  3.620 2.700 3.860 3.400 ;
        RECT  0.560 2.700 0.780 3.880 ;
        RECT  3.700 2.700 3.860 4.180 ;
        RECT  3.700 3.910 3.980 4.180 ;
        RECT  0.770 0.300 4.440 0.460 ;
        RECT  4.140 0.300 4.440 0.570 ;
        RECT  0.770 0.300 0.930 0.860 ;
        RECT  0.470 0.580 0.930 0.860 ;
        RECT  0.420 1.690 0.660 2.100 ;
        RECT  4.200 1.890 4.540 2.100 ;
        RECT  0.420 1.940 4.540 2.100 ;
        RECT  4.440 3.020 4.940 3.260 ;
        RECT  2.280 3.450 2.480 4.100 ;
        RECT  2.280 3.940 3.540 4.100 ;
        RECT  3.380 3.940 3.540 4.500 ;
        RECT  4.260 3.980 4.600 4.500 ;
        RECT  4.440 3.020 4.600 4.500 ;
        RECT  3.380 4.340 4.600 4.500 ;
        RECT  4.050 1.070 5.770 1.230 ;
        RECT  4.050 1.070 4.340 1.390 ;
        RECT  5.570 0.620 5.770 1.780 ;
        RECT  5.570 1.620 5.970 1.780 ;
        RECT  5.650 3.020 7.170 3.220 ;
        RECT  6.890 3.020 7.170 3.460 ;
        RECT  5.650 3.020 5.810 4.180 ;
        RECT  5.430 3.880 5.810 4.180 ;
        RECT  3.290 1.550 4.860 1.710 ;
        RECT  3.290 1.550 3.650 1.780 ;
        RECT  4.700 1.550 4.860 2.100 ;
        RECT  4.700 1.940 7.680 2.100 ;
        RECT  6.010 3.940 7.820 4.100 ;
        RECT  4.760 3.420 4.920 4.500 ;
        RECT  6.010 3.940 6.170 4.500 ;
        RECT  4.760 4.340 6.170 4.500 ;
        RECT  6.970 0.640 7.250 1.240 ;
        RECT  6.970 0.960 7.850 1.240 ;
        RECT  6.970 0.640 7.130 1.760 ;
        RECT  6.710 1.500 7.130 1.760 ;
        RECT  5.990 3.500 6.290 3.780 ;
        RECT  5.990 3.620 8.630 3.780 ;
        RECT  8.350 3.340 8.630 4.420 ;
        RECT  8.180 3.620 8.630 4.420 ;
        RECT  4.120 2.700 8.940 2.860 ;
        RECT  5.220 2.700 5.420 3.690 ;
        RECT  4.120 2.700 4.280 3.740 ;
        RECT  4.020 3.340 4.280 3.740 ;
        RECT  7.330 3.020 9.170 3.180 ;
        RECT  7.330 3.020 7.530 3.310 ;
        RECT  8.970 3.020 9.170 3.380 ;
        RECT  5.090 0.300 6.100 0.460 ;
        RECT  6.580 0.300 8.890 0.460 ;
        RECT  5.940 0.300 6.100 0.740 ;
        RECT  8.730 0.300 8.890 0.740 ;
        RECT  6.580 0.300 6.740 0.740 ;
        RECT  5.940 0.580 6.740 0.740 ;
        RECT  8.730 0.580 9.170 0.740 ;
        RECT  3.080 0.620 3.980 0.780 ;
        RECT  5.090 0.300 5.330 0.910 ;
        RECT  3.820 0.750 5.330 0.910 ;
        RECT  7.910 0.620 8.250 0.780 ;
        RECT  8.010 0.620 8.250 1.410 ;
        RECT  8.010 1.250 9.230 1.410 ;
        RECT  8.920 1.250 9.230 1.690 ;
        RECT  8.010 0.620 8.190 1.710 ;
        RECT  7.460 1.490 8.190 1.710 ;
        RECT  9.160 3.570 9.320 4.380 ;
        RECT  8.920 4.220 9.320 4.380 ;
        LAYER VTPH ;
        RECT  0.000 1.160 1.130 3.660 ;
        RECT  2.980 1.210 4.190 3.540 ;
        RECT  6.020 1.160 9.600 3.540 ;
        RECT  0.000 1.260 9.600 3.540 ;
        RECT  0.000 1.260 4.120 3.600 ;
        RECT  0.000 1.260 2.810 3.660 ;
        RECT  8.380 1.140 9.600 3.660 ;
        RECT  7.030 1.160 9.060 3.860 ;
        LAYER VTNH ;
        RECT  2.810 3.600 7.030 4.800 ;
        RECT  4.120 3.540 7.030 4.800 ;
        RECT  0.000 3.660 7.030 4.800 ;
        RECT  9.060 3.660 9.600 4.800 ;
        RECT  0.000 3.860 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  0.000 0.000 8.380 1.160 ;
        RECT  1.130 0.000 6.020 1.210 ;
        RECT  1.130 0.000 2.980 1.260 ;
        RECT  4.190 0.000 6.020 1.260 ;
    END
END SDFERM1HM

MACRO SDFEQZRM8HM
    CLASS CORE ;
    FOREIGN SDFEQZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.047  LAYER ME1  ;
        ANTENNAGATEAREA 0.047  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.222  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 3.500 1.100 3.700 ;
        LAYER ME2 ;
        RECT  0.900 3.420 1.100 3.960 ;
        LAYER ME1 ;
        RECT  0.860 3.380 1.260 3.810 ;
        END
    END SD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        ANTENNAGATEAREA 0.140  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.630  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.150 5.100 1.350 ;
        LAYER ME2 ;
        RECT  4.900 1.090 5.100 1.970 ;
        LAYER ME1 ;
        RECT  4.560 1.030 5.200 1.370 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 3.400 3.600 3.900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.840 1.600 1.330 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.800 0.780 1.330 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.007  LAYER ME1  ;
        ANTENNADIFFAREA 0.965  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.250 2.730 9.530 4.450 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 3.490 2.560 3.680 ;
        RECT  0.540 3.970 1.900 4.130 ;
        RECT  1.500 3.490 1.900 4.130 ;
        RECT  0.480 3.690 0.700 3.970 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.830 1.610 9.990 2.910 ;
        RECT  8.750 1.580 8.970 2.860 ;
        RECT  7.330 2.260 7.530 3.500 ;
        RECT  2.510 2.180 2.790 2.540 ;
        RECT  0.750 2.260 1.030 2.860 ;
        RECT  0.680 1.810 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.830 -0.140 9.990 0.750 ;
        RECT  8.730 -0.140 8.990 0.710 ;
        RECT  7.690 -0.140 7.850 0.750 ;
        RECT  4.420 -0.140 4.700 0.530 ;
        RECT  0.700 -0.140 0.960 0.640 ;
        RECT  0.000 4.660 10.400 4.940 ;
        RECT  9.780 4.170 9.990 4.940 ;
        RECT  8.770 4.170 8.990 4.940 ;
        RECT  7.300 4.200 7.530 4.940 ;
        RECT  5.070 4.480 5.350 4.940 ;
        RECT  3.070 4.480 3.350 4.940 ;
        RECT  0.740 4.300 1.020 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.470 2.810 1.750 3.180 ;
        RECT  0.140 3.020 1.750 3.180 ;
        RECT  0.140 3.020 0.360 3.340 ;
        RECT  0.140 3.020 0.300 4.500 ;
        RECT  0.140 4.240 0.420 4.500 ;
        RECT  0.100 0.390 0.380 0.650 ;
        RECT  1.810 0.980 2.510 1.260 ;
        RECT  0.100 0.390 0.300 1.970 ;
        RECT  0.940 1.070 1.100 1.650 ;
        RECT  1.810 0.980 1.970 1.650 ;
        RECT  0.100 1.490 1.970 1.650 ;
        RECT  0.100 1.490 0.420 1.970 ;
        RECT  2.500 3.060 3.060 3.220 ;
        RECT  2.900 3.060 3.060 4.000 ;
        RECT  2.310 3.840 3.060 4.000 ;
        RECT  2.310 3.840 2.590 4.180 ;
        RECT  2.120 0.620 3.430 0.780 ;
        RECT  3.270 0.620 3.430 1.460 ;
        RECT  2.720 1.300 3.430 1.460 ;
        RECT  2.720 1.300 2.880 1.630 ;
        RECT  2.600 1.470 2.760 2.020 ;
        RECT  1.540 1.860 2.760 2.020 ;
        RECT  3.620 0.620 3.920 0.870 ;
        RECT  3.620 0.620 3.860 1.780 ;
        RECT  3.040 1.620 3.860 1.780 ;
        RECT  3.040 1.620 3.200 2.070 ;
        RECT  2.920 1.850 3.200 2.070 ;
        RECT  3.620 3.020 4.110 3.180 ;
        RECT  3.830 3.020 4.110 4.180 ;
        RECT  4.070 1.020 4.350 1.760 ;
        RECT  4.070 1.600 5.100 1.760 ;
        RECT  1.180 0.300 4.260 0.460 ;
        RECT  1.180 0.300 1.460 0.610 ;
        RECT  4.100 0.300 4.260 0.850 ;
        RECT  5.000 0.380 5.160 0.850 ;
        RECT  4.100 0.690 5.160 0.850 ;
        RECT  1.930 2.700 5.670 2.860 ;
        RECT  1.930 2.700 2.150 3.320 ;
        RECT  5.550 4.080 5.830 4.290 ;
        RECT  4.750 4.130 5.830 4.290 ;
        RECT  2.750 4.160 3.670 4.320 ;
        RECT  3.510 4.160 3.670 4.500 ;
        RECT  2.750 4.160 2.910 4.500 ;
        RECT  1.640 4.340 2.910 4.500 ;
        RECT  4.750 4.130 4.910 4.500 ;
        RECT  3.510 4.340 4.910 4.500 ;
        RECT  4.740 3.020 5.020 3.360 ;
        RECT  4.740 3.200 6.710 3.360 ;
        RECT  4.740 3.020 4.960 3.560 ;
        RECT  4.310 3.400 4.960 3.560 ;
        RECT  6.550 3.200 6.710 4.130 ;
        RECT  4.310 3.400 4.590 4.180 ;
        RECT  6.570 2.720 6.850 2.970 ;
        RECT  5.830 2.810 7.090 2.970 ;
        RECT  6.930 2.810 7.090 4.460 ;
        RECT  6.130 4.300 7.090 4.460 ;
        RECT  6.860 0.660 7.140 1.680 ;
        RECT  6.860 1.430 7.760 1.680 ;
        RECT  6.580 1.530 7.050 1.780 ;
        RECT  6.060 0.340 7.530 0.500 ;
        RECT  7.370 0.340 7.530 1.230 ;
        RECT  7.370 0.950 7.950 1.230 ;
        RECT  6.060 0.340 6.340 1.730 ;
        RECT  7.880 2.730 8.240 4.500 ;
        RECT  5.420 0.340 5.700 0.630 ;
        RECT  5.470 0.340 5.700 2.100 ;
        RECT  3.360 1.940 8.280 2.100 ;
        RECT  8.200 0.400 8.520 1.280 ;
        RECT  8.200 0.990 9.080 1.280 ;
        RECT  8.200 0.400 8.440 1.770 ;
        RECT  8.070 1.490 8.440 1.770 ;
        RECT  9.310 0.400 9.540 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.620 3.660 ;
        RECT  7.310 1.140 10.400 3.660 ;
        RECT  5.550 1.180 8.420 3.710 ;
        RECT  6.970 1.180 8.420 3.900 ;
        LAYER VTNH ;
        RECT  0.000 3.660 5.550 4.800 ;
        RECT  0.000 3.710 6.970 4.800 ;
        RECT  8.420 3.660 10.400 4.800 ;
        RECT  0.000 3.900 10.400 4.800 ;
        RECT  0.000 0.000 10.400 1.140 ;
        RECT  6.620 0.000 7.310 1.180 ;
    END
END SDFEQZRM8HM

MACRO SDFEQZRM4HM
    CLASS CORE ;
    FOREIGN SDFEQZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.992  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 3.500 1.100 3.700 ;
        LAYER ME2 ;
        RECT  0.900 3.420 1.100 3.960 ;
        LAYER ME1 ;
        RECT  0.860 3.380 1.260 3.810 ;
        END
    END SD
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        ANTENNAGATEAREA 0.148  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.629  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.150 5.100 1.350 ;
        LAYER ME2 ;
        RECT  4.900 1.090 5.100 1.970 ;
        LAYER ME1 ;
        RECT  4.560 1.030 5.250 1.370 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 3.400 3.600 3.900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.840 1.700 1.330 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.800 0.780 1.330 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.018  LAYER ME1  ;
        ANTENNADIFFAREA 0.841  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.190 2.730 9.500 4.450 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 3.490 2.560 3.680 ;
        RECT  0.540 3.970 2.000 4.130 ;
        RECT  1.500 3.490 2.000 4.130 ;
        RECT  0.480 3.690 0.700 3.970 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.690 1.660 8.910 2.950 ;
        RECT  7.330 2.260 7.530 3.500 ;
        RECT  2.510 2.180 2.790 2.540 ;
        RECT  0.750 2.260 1.030 2.860 ;
        RECT  0.680 1.810 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.670 -0.140 8.930 0.710 ;
        RECT  7.690 -0.140 7.850 0.750 ;
        RECT  4.420 -0.140 4.700 0.530 ;
        RECT  0.700 -0.140 0.960 0.640 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  8.710 4.170 8.930 4.940 ;
        RECT  7.300 4.200 7.530 4.940 ;
        RECT  5.070 4.480 5.350 4.940 ;
        RECT  3.070 4.480 3.350 4.940 ;
        RECT  0.740 4.300 1.020 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.470 2.810 1.750 3.180 ;
        RECT  0.140 3.020 1.750 3.180 ;
        RECT  0.140 3.020 0.360 3.340 ;
        RECT  0.140 3.020 0.300 4.500 ;
        RECT  0.140 4.240 0.420 4.500 ;
        RECT  0.100 0.390 0.380 0.650 ;
        RECT  2.030 0.980 2.510 1.260 ;
        RECT  0.100 0.390 0.300 1.970 ;
        RECT  0.940 1.070 1.100 1.650 ;
        RECT  2.030 0.980 2.190 1.650 ;
        RECT  0.100 1.490 2.190 1.650 ;
        RECT  0.100 1.490 0.420 1.970 ;
        RECT  2.500 3.060 3.060 3.220 ;
        RECT  2.900 3.060 3.060 4.000 ;
        RECT  2.310 3.840 3.060 4.000 ;
        RECT  2.310 3.840 2.590 4.180 ;
        RECT  2.120 0.620 3.430 0.780 ;
        RECT  3.270 0.620 3.430 1.460 ;
        RECT  2.720 1.300 3.430 1.460 ;
        RECT  2.720 1.300 2.880 1.630 ;
        RECT  2.600 1.470 2.760 2.020 ;
        RECT  1.540 1.860 2.760 2.020 ;
        RECT  3.620 0.620 3.920 0.870 ;
        RECT  3.620 0.620 3.860 1.780 ;
        RECT  3.040 1.620 3.860 1.780 ;
        RECT  3.040 1.620 3.200 2.070 ;
        RECT  2.920 1.850 3.200 2.070 ;
        RECT  3.620 3.070 4.110 3.230 ;
        RECT  3.830 3.070 4.110 4.180 ;
        RECT  4.070 1.020 4.350 1.760 ;
        RECT  4.070 1.600 5.100 1.760 ;
        RECT  1.180 0.300 4.260 0.460 ;
        RECT  1.180 0.300 1.460 0.610 ;
        RECT  4.100 0.300 4.260 0.850 ;
        RECT  5.000 0.380 5.160 0.850 ;
        RECT  4.100 0.690 5.160 0.850 ;
        RECT  1.930 2.700 5.670 2.860 ;
        RECT  1.930 2.700 2.150 3.320 ;
        RECT  5.550 4.080 5.830 4.290 ;
        RECT  4.750 4.130 5.830 4.290 ;
        RECT  2.750 4.160 3.670 4.320 ;
        RECT  3.510 4.160 3.670 4.500 ;
        RECT  2.750 4.160 2.910 4.500 ;
        RECT  1.640 4.340 2.910 4.500 ;
        RECT  4.750 4.130 4.910 4.500 ;
        RECT  3.510 4.340 4.910 4.500 ;
        RECT  4.740 3.020 5.020 3.360 ;
        RECT  4.740 3.200 6.710 3.360 ;
        RECT  4.740 3.020 4.960 3.560 ;
        RECT  4.310 3.400 4.960 3.560 ;
        RECT  6.550 3.200 6.710 4.130 ;
        RECT  4.310 3.400 4.590 4.180 ;
        RECT  6.570 2.720 6.850 2.970 ;
        RECT  5.830 2.810 7.090 2.970 ;
        RECT  6.930 2.810 7.090 4.460 ;
        RECT  6.130 4.300 7.090 4.460 ;
        RECT  6.860 0.660 7.140 1.680 ;
        RECT  6.860 1.430 7.760 1.680 ;
        RECT  6.580 1.530 7.050 1.780 ;
        RECT  6.060 0.340 7.530 0.500 ;
        RECT  7.370 0.340 7.530 1.230 ;
        RECT  7.370 0.950 7.950 1.230 ;
        RECT  6.060 0.340 6.340 1.730 ;
        RECT  7.880 2.730 8.180 4.500 ;
        RECT  5.420 0.340 5.700 0.630 ;
        RECT  5.470 0.340 5.700 2.100 ;
        RECT  3.360 1.940 8.220 2.100 ;
        RECT  8.140 0.400 8.460 1.280 ;
        RECT  8.140 0.990 9.020 1.280 ;
        RECT  8.140 0.400 8.330 1.770 ;
        RECT  8.010 1.490 8.330 1.770 ;
        RECT  9.250 0.400 9.470 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.620 3.660 ;
        RECT  7.310 1.140 9.600 3.660 ;
        RECT  5.550 1.180 8.420 3.710 ;
        RECT  6.970 1.180 8.420 3.800 ;
        LAYER VTNH ;
        RECT  0.000 3.660 5.550 4.800 ;
        RECT  0.000 3.710 6.970 4.800 ;
        RECT  8.420 3.660 9.600 4.800 ;
        RECT  0.000 3.800 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  6.620 0.000 7.310 1.180 ;
    END
END SDFEQZRM4HM

MACRO SDFEQZRM2HM
    CLASS CORE ;
    FOREIGN SDFEQZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        ANTENNAGATEAREA 0.148  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.629  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.150 5.100 1.350 ;
        LAYER ME2 ;
        RECT  4.900 1.090 5.100 1.970 ;
        LAYER ME1 ;
        RECT  4.560 1.030 5.250 1.370 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.992  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 3.500 1.100 3.700 ;
        LAYER ME2 ;
        RECT  0.900 3.420 1.100 3.960 ;
        LAYER ME1 ;
        RECT  0.860 3.380 1.260 3.810 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 3.400 3.600 3.900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.840 1.700 1.330 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.800 0.780 1.330 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.070 2.780 9.350 4.450 ;
        RECT  8.840 3.240 9.350 3.560 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 3.490 2.560 3.680 ;
        RECT  0.540 3.970 2.000 4.130 ;
        RECT  1.500 3.490 2.000 4.130 ;
        RECT  0.480 3.690 0.700 3.970 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.690 1.660 8.910 2.540 ;
        RECT  8.570 2.260 8.790 3.000 ;
        RECT  7.330 2.260 7.530 3.500 ;
        RECT  2.510 2.180 2.790 2.540 ;
        RECT  0.750 2.260 1.030 2.860 ;
        RECT  0.680 1.810 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.670 -0.140 8.940 0.710 ;
        RECT  7.690 -0.140 7.850 0.750 ;
        RECT  4.420 -0.140 4.700 0.530 ;
        RECT  0.700 -0.140 0.960 0.640 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  8.590 4.170 8.810 4.940 ;
        RECT  7.300 4.200 7.530 4.940 ;
        RECT  5.070 4.480 5.350 4.940 ;
        RECT  3.070 4.480 3.350 4.940 ;
        RECT  0.740 4.300 1.020 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.470 2.810 1.750 3.180 ;
        RECT  0.140 3.020 1.750 3.180 ;
        RECT  0.140 3.020 0.360 3.340 ;
        RECT  0.140 3.020 0.300 4.500 ;
        RECT  0.140 4.240 0.420 4.500 ;
        RECT  0.100 0.390 0.380 0.650 ;
        RECT  2.030 0.980 2.510 1.260 ;
        RECT  0.100 0.390 0.300 1.970 ;
        RECT  0.940 1.070 1.100 1.650 ;
        RECT  2.030 0.980 2.190 1.650 ;
        RECT  0.100 1.490 2.190 1.650 ;
        RECT  0.100 1.490 0.420 1.970 ;
        RECT  2.500 3.060 3.060 3.220 ;
        RECT  2.900 3.060 3.060 4.000 ;
        RECT  2.310 3.840 3.060 4.000 ;
        RECT  2.310 3.840 2.590 4.180 ;
        RECT  2.120 0.620 3.430 0.780 ;
        RECT  3.270 0.620 3.430 1.460 ;
        RECT  2.720 1.300 3.430 1.460 ;
        RECT  2.720 1.300 2.880 1.630 ;
        RECT  2.600 1.470 2.760 2.020 ;
        RECT  1.540 1.860 2.760 2.020 ;
        RECT  3.620 0.620 3.920 0.870 ;
        RECT  3.620 0.620 3.860 1.780 ;
        RECT  3.040 1.620 3.860 1.780 ;
        RECT  3.040 1.620 3.200 2.070 ;
        RECT  2.920 1.850 3.200 2.070 ;
        RECT  3.620 3.070 4.110 3.230 ;
        RECT  3.830 3.070 4.110 4.180 ;
        RECT  4.070 1.020 4.350 1.760 ;
        RECT  4.070 1.600 5.100 1.760 ;
        RECT  1.180 0.300 4.260 0.460 ;
        RECT  1.180 0.300 1.460 0.610 ;
        RECT  4.100 0.300 4.260 0.850 ;
        RECT  5.000 0.380 5.160 0.850 ;
        RECT  4.100 0.690 5.160 0.850 ;
        RECT  1.930 2.700 5.670 2.860 ;
        RECT  1.930 2.700 2.150 3.320 ;
        RECT  5.550 4.080 5.830 4.290 ;
        RECT  4.750 4.130 5.830 4.290 ;
        RECT  2.750 4.160 3.670 4.320 ;
        RECT  3.510 4.160 3.670 4.500 ;
        RECT  2.750 4.160 2.910 4.500 ;
        RECT  1.640 4.340 2.910 4.500 ;
        RECT  4.750 4.130 4.910 4.500 ;
        RECT  3.510 4.340 4.910 4.500 ;
        RECT  4.740 3.020 5.020 3.360 ;
        RECT  4.740 3.200 6.710 3.360 ;
        RECT  4.740 3.020 4.960 3.560 ;
        RECT  4.310 3.400 4.960 3.560 ;
        RECT  6.550 3.200 6.710 4.130 ;
        RECT  4.310 3.400 4.590 4.180 ;
        RECT  6.570 2.720 6.850 2.970 ;
        RECT  5.830 2.810 7.090 2.970 ;
        RECT  6.930 2.810 7.090 4.460 ;
        RECT  6.130 4.300 7.090 4.460 ;
        RECT  6.860 0.660 7.140 1.680 ;
        RECT  6.860 1.430 7.760 1.680 ;
        RECT  6.580 1.530 7.050 1.780 ;
        RECT  6.060 0.340 7.530 0.500 ;
        RECT  7.370 0.340 7.530 1.230 ;
        RECT  7.370 0.950 7.950 1.230 ;
        RECT  6.060 0.340 6.340 1.730 ;
        RECT  7.880 2.730 8.180 4.500 ;
        RECT  5.420 0.340 5.700 0.630 ;
        RECT  5.470 0.340 5.700 2.100 ;
        RECT  3.360 1.940 8.220 2.100 ;
        RECT  8.140 0.400 8.460 1.280 ;
        RECT  8.140 0.990 9.020 1.280 ;
        RECT  8.140 0.400 8.330 1.770 ;
        RECT  8.010 1.490 8.330 1.770 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.620 3.660 ;
        RECT  7.310 1.140 9.600 3.660 ;
        RECT  5.550 1.180 8.420 3.710 ;
        RECT  6.970 1.180 8.420 3.800 ;
        LAYER VTNH ;
        RECT  0.000 3.660 5.550 4.800 ;
        RECT  0.000 3.710 6.970 4.800 ;
        RECT  8.420 3.660 9.600 4.800 ;
        RECT  0.000 3.800 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  6.620 0.000 7.310 1.180 ;
    END
END SDFEQZRM2HM

MACRO SDFEQZRM1HM
    CLASS CORE ;
    FOREIGN SDFEQZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.068  LAYER ME1  ;
        ANTENNAGATEAREA 0.068  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.538  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.230 3.900 1.430 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.480 1.160 4.070 1.430 ;
        END
    END SD
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.470 3.620 5.910 4.070 ;
        RECT  5.670 3.530 5.910 4.070 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 3.600 2.480 4.000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.670 3.520 1.900 3.990 ;
        RECT  0.420 3.520 1.900 3.680 ;
        RECT  0.420 3.520 0.640 3.810 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.112  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.180 3.940 8.450 4.310 ;
        RECT  8.210 2.980 8.450 4.310 ;
        RECT  7.230 3.940 8.450 4.100 ;
        RECT  7.230 3.550 7.570 4.100 ;
        RECT  3.990 4.340 7.450 4.500 ;
        RECT  7.230 3.550 7.450 4.500 ;
        RECT  3.990 3.320 4.150 4.500 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 3.840 1.240 4.300 ;
        END
    END RB
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.750 1.200 0.970 ;
        RECT  0.500 0.750 0.770 1.160 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.630 2.260 7.910 2.810 ;
        RECT  5.550 2.260 5.840 2.580 ;
        RECT  4.110 2.260 4.390 3.020 ;
        RECT  2.390 2.260 2.670 2.720 ;
        RECT  0.820 1.930 1.100 2.540 ;
        RECT  0.620 2.260 0.900 3.000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  6.610 -0.140 6.890 0.500 ;
        RECT  2.640 -0.140 2.920 0.320 ;
        RECT  0.660 -0.140 0.940 0.580 ;
        RECT  0.000 4.660 8.800 4.940 ;
        RECT  7.610 4.400 7.890 4.940 ;
        RECT  0.730 4.480 1.010 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.000 1.160 2.760 1.320 ;
        RECT  1.000 1.160 1.160 1.770 ;
        RECT  0.100 1.610 1.160 1.770 ;
        RECT  0.100 0.330 0.340 1.880 ;
        RECT  1.140 0.300 2.470 0.460 ;
        RECT  2.300 0.300 2.470 0.680 ;
        RECT  1.140 0.300 1.450 0.570 ;
        RECT  2.300 0.520 3.580 0.680 ;
        RECT  1.180 2.730 2.040 3.040 ;
        RECT  1.180 2.880 3.590 3.040 ;
        RECT  3.130 2.880 3.290 4.180 ;
        RECT  2.980 3.950 3.290 4.180 ;
        RECT  0.100 2.780 0.380 3.360 ;
        RECT  0.100 3.200 2.900 3.360 ;
        RECT  2.640 3.200 2.900 3.590 ;
        RECT  0.100 2.780 0.260 4.440 ;
        RECT  2.640 3.200 2.820 4.500 ;
        RECT  0.100 4.150 0.380 4.440 ;
        RECT  3.480 3.510 3.640 4.500 ;
        RECT  2.640 4.340 3.640 4.500 ;
        RECT  4.230 0.620 4.540 0.840 ;
        RECT  3.010 1.160 3.290 1.750 ;
        RECT  4.230 0.620 4.410 1.750 ;
        RECT  3.010 1.590 4.410 1.750 ;
        RECT  1.740 1.640 2.420 2.100 ;
        RECT  4.560 1.820 4.910 2.100 ;
        RECT  1.740 1.940 4.910 2.100 ;
        RECT  3.770 0.300 5.130 0.460 ;
        RECT  4.850 0.300 5.130 0.500 ;
        RECT  1.720 0.620 2.000 1.000 ;
        RECT  3.770 0.300 3.930 1.000 ;
        RECT  1.720 0.840 3.930 1.000 ;
        RECT  5.130 3.060 6.340 3.260 ;
        RECT  5.130 3.060 5.520 3.420 ;
        RECT  6.070 3.060 6.340 4.130 ;
        RECT  6.070 3.470 6.570 3.760 ;
        RECT  6.070 3.470 6.350 4.130 ;
        RECT  5.530 0.330 5.810 1.140 ;
        RECT  5.390 0.980 7.080 1.140 ;
        RECT  5.390 0.960 5.590 1.750 ;
        RECT  6.040 2.700 7.220 2.860 ;
        RECT  4.650 2.740 6.200 2.900 ;
        RECT  4.650 2.740 4.880 4.130 ;
        RECT  4.650 3.910 5.240 4.130 ;
        RECT  7.130 0.340 7.460 0.820 ;
        RECT  6.160 0.660 7.460 0.820 ;
        RECT  6.210 1.620 7.980 1.780 ;
        RECT  6.500 3.050 8.050 3.230 ;
        RECT  6.500 3.050 6.920 3.260 ;
        RECT  7.770 3.050 8.050 3.760 ;
        RECT  6.760 3.050 6.920 4.180 ;
        RECT  6.560 3.950 6.920 4.180 ;
        RECT  4.860 0.750 5.230 1.050 ;
        RECT  7.820 1.030 8.100 1.460 ;
        RECT  5.830 1.300 8.100 1.460 ;
        RECT  5.070 0.750 5.230 2.070 ;
        RECT  5.830 1.300 5.990 2.070 ;
        RECT  5.070 1.910 5.990 2.070 ;
        RECT  7.720 0.340 8.530 0.500 ;
        RECT  8.370 0.340 8.530 1.970 ;
        RECT  8.230 1.680 8.530 1.970 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 3.540 ;
        RECT  5.130 1.140 8.800 3.600 ;
        RECT  0.000 1.140 2.530 3.660 ;
        RECT  6.800 1.140 8.800 3.660 ;
        LAYER VTNH ;
        RECT  2.530 3.540 5.130 4.800 ;
        RECT  2.530 3.600 6.800 4.800 ;
        RECT  0.000 3.660 8.800 4.800 ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END SDFEQZRM1HM

MACRO SDFEQRM8HM
    CLASS CORE ;
    FOREIGN SDFEQRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.108  LAYER ME1  ;
        ANTENNAGATEAREA 0.108  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.659  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.050 1.070 4.250 1.270 ;
        LAYER ME2 ;
        RECT  4.010 0.840 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.920 0.950 4.280 1.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.901  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.170 1.050 7.370 1.250 ;
        LAYER ME2 ;
        RECT  7.170 0.840 7.500 1.560 ;
        LAYER ME1 ;
        RECT  7.000 0.900 7.370 1.340 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 3.370  LAYER ME1  ;
        ANTENNADIFFAREA 1.417  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 2.900 1.640 3.100 ;
        RECT  1.440 3.960 1.600 4.390 ;
        RECT  0.100 3.960 1.600 4.120 ;
        RECT  0.100 2.900 0.340 4.460 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        ANTENNAGATEAREA 0.199  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.141  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.560 1.110 6.760 1.310 ;
        LAYER ME2 ;
        RECT  6.500 0.840 6.760 1.560 ;
        LAYER ME1 ;
        RECT  6.560 0.900 6.820 1.460 ;
        END
    END E
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.293  LAYER ME1  ;
        ANTENNAGATEAREA 0.293  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.458  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 3.550 3.500 3.750 ;
        LAYER ME2 ;
        RECT  3.300 3.240 3.500 3.960 ;
        LAYER ME1 ;
        RECT  3.240 3.540 3.940 3.750 ;
        RECT  3.240 3.340 3.560 3.750 ;
        RECT  2.130 3.340 3.560 3.500 ;
        RECT  2.130 3.340 2.290 3.790 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.425  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 0.780 3.100 0.980 ;
        LAYER ME2 ;
        RECT  2.900 0.440 3.100 1.160 ;
        LAYER ME1 ;
        RECT  2.740 0.710 3.280 1.040 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.163  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.460 1.100 3.660 1.300 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.660 1.560 ;
        LAYER ME1 ;
        RECT  2.170 1.200 3.760 1.360 ;
        RECT  3.460 1.030 3.760 1.360 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.220 1.570 9.510 2.540 ;
        RECT  0.680 1.780 0.970 2.720 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  6.890 -0.140 7.050 0.420 ;
        RECT  0.660 -0.140 0.940 0.380 ;
        RECT  0.000 4.660 10.400 4.940 ;
        RECT  7.130 4.260 7.410 4.940 ;
        RECT  3.800 4.260 4.080 4.940 ;
        RECT  1.900 4.270 2.180 4.940 ;
        RECT  0.620 4.280 0.900 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.390 0.320 2.020 ;
        RECT  1.680 0.740 2.460 0.900 ;
        RECT  1.030 1.080 1.840 1.240 ;
        RECT  1.680 0.740 1.840 1.780 ;
        RECT  1.680 1.550 3.760 1.780 ;
        RECT  1.800 3.020 4.320 3.180 ;
        RECT  0.600 3.570 1.970 3.730 ;
        RECT  4.160 3.020 4.320 3.740 ;
        RECT  1.800 3.020 1.970 4.110 ;
        RECT  1.800 3.950 2.500 4.110 ;
        RECT  2.340 3.950 2.500 4.450 ;
        RECT  2.340 4.290 3.160 4.450 ;
        RECT  4.480 2.700 4.790 2.920 ;
        RECT  4.480 2.700 4.720 3.400 ;
        RECT  4.560 2.700 4.720 4.180 ;
        RECT  4.560 3.910 4.840 4.180 ;
        RECT  1.360 0.300 5.070 0.460 ;
        RECT  4.770 0.300 5.070 0.570 ;
        RECT  1.360 0.300 1.520 0.800 ;
        RECT  1.160 0.640 1.520 0.800 ;
        RECT  1.260 1.780 1.500 2.100 ;
        RECT  4.830 1.890 5.170 2.100 ;
        RECT  1.260 1.940 5.170 2.100 ;
        RECT  5.300 3.020 5.800 3.260 ;
        RECT  2.660 3.660 2.940 4.100 ;
        RECT  2.660 3.940 4.400 4.100 ;
        RECT  4.240 3.940 4.400 4.500 ;
        RECT  5.120 3.980 5.460 4.500 ;
        RECT  5.300 3.020 5.460 4.500 ;
        RECT  4.240 4.340 5.460 4.500 ;
        RECT  4.680 1.070 6.400 1.230 ;
        RECT  4.680 1.070 4.970 1.390 ;
        RECT  6.200 0.620 6.400 1.780 ;
        RECT  6.200 1.620 6.600 1.780 ;
        RECT  6.450 3.020 7.970 3.220 ;
        RECT  7.690 3.020 7.970 3.460 ;
        RECT  6.450 3.020 6.610 4.180 ;
        RECT  6.020 3.850 6.610 4.180 ;
        RECT  3.920 1.550 5.490 1.710 ;
        RECT  3.920 1.550 4.280 1.780 ;
        RECT  5.330 1.550 5.490 2.100 ;
        RECT  5.330 1.940 8.090 2.100 ;
        RECT  6.810 3.940 8.620 4.100 ;
        RECT  5.620 3.420 5.780 4.500 ;
        RECT  6.810 3.940 6.970 4.500 ;
        RECT  5.620 4.340 6.970 4.500 ;
        RECT  7.530 0.640 7.810 1.180 ;
        RECT  7.530 1.020 8.710 1.180 ;
        RECT  7.530 0.640 7.690 1.760 ;
        RECT  7.270 1.500 7.690 1.760 ;
        RECT  6.790 3.500 7.090 3.780 ;
        RECT  6.790 3.620 9.430 3.780 ;
        RECT  9.150 3.340 9.430 4.420 ;
        RECT  8.980 3.620 9.430 4.420 ;
        RECT  5.720 0.300 6.730 0.460 ;
        RECT  7.210 0.300 9.400 0.460 ;
        RECT  6.570 0.300 6.730 0.740 ;
        RECT  9.240 0.300 9.400 0.740 ;
        RECT  7.210 0.300 7.370 0.740 ;
        RECT  6.570 0.580 7.370 0.740 ;
        RECT  9.240 0.580 9.680 0.740 ;
        RECT  3.710 0.620 4.610 0.780 ;
        RECT  5.720 0.300 5.960 0.910 ;
        RECT  4.450 0.750 5.960 0.910 ;
        RECT  4.980 2.700 9.740 2.860 ;
        RECT  6.080 2.700 6.280 3.670 ;
        RECT  4.980 2.700 5.140 3.740 ;
        RECT  4.880 3.340 5.140 3.740 ;
        RECT  8.130 3.020 9.970 3.180 ;
        RECT  8.130 3.020 8.330 3.310 ;
        RECT  9.770 3.020 9.970 3.380 ;
        RECT  8.490 0.620 9.060 0.780 ;
        RECT  8.900 1.250 10.030 1.410 ;
        RECT  8.900 0.620 9.060 1.680 ;
        RECT  7.870 1.460 9.060 1.680 ;
        RECT  9.720 1.250 10.030 1.690 ;
        RECT  9.960 3.570 10.120 4.380 ;
        RECT  9.720 4.220 10.120 4.380 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.010 3.660 ;
        RECT  3.610 1.210 4.820 3.600 ;
        RECT  6.650 1.160 10.400 3.540 ;
        RECT  0.000 1.260 10.400 3.540 ;
        RECT  0.000 1.260 4.980 3.600 ;
        RECT  0.000 1.260 3.670 3.660 ;
        RECT  9.070 1.140 10.400 3.660 ;
        RECT  7.830 1.160 9.860 3.860 ;
        LAYER VTNH ;
        RECT  3.670 3.600 7.830 4.800 ;
        RECT  4.980 3.540 7.830 4.800 ;
        RECT  0.000 3.660 7.830 4.800 ;
        RECT  9.860 3.660 10.400 4.800 ;
        RECT  0.000 3.860 10.400 4.800 ;
        RECT  0.000 0.000 10.400 1.140 ;
        RECT  1.010 0.000 9.070 1.160 ;
        RECT  1.010 0.000 6.650 1.210 ;
        RECT  1.010 0.000 3.610 1.260 ;
        RECT  4.820 0.000 6.650 1.260 ;
    END
END SDFEQRM8HM

MACRO SDFEQRM4HM
    CLASS CORE ;
    FOREIGN SDFEQRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.985  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.850 3.550 3.050 3.750 ;
        LAYER ME2 ;
        RECT  2.850 3.240 3.100 3.960 ;
        LAYER ME1 ;
        RECT  2.620 3.340 3.140 3.750 ;
        END
    END RB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        ANTENNAGATEAREA 0.199  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.141  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.930 1.110 6.130 1.310 ;
        LAYER ME2 ;
        RECT  5.700 0.840 6.130 1.560 ;
        LAYER ME1 ;
        RECT  5.930 0.900 6.190 1.460 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        ANTENNAGATEAREA 0.118  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.361  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.070 3.500 1.270 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.290 0.950 3.650 1.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.370 0.900 6.810 1.340 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.498  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 3.040 1.100 4.390 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        ANTENNAGATEAREA 0.048  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.183  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 0.780 2.300 0.980 ;
        LAYER ME2 ;
        RECT  2.100 0.440 2.300 1.160 ;
        LAYER ME1 ;
        RECT  2.040 0.710 2.650 1.040 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER ME1  ;
        ANTENNAGATEAREA 0.162  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.163  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.100 3.100 1.300 ;
        LAYER ME2 ;
        RECT  2.900 0.840 3.100 1.560 ;
        LAYER ME1 ;
        RECT  1.540 1.200 3.130 1.360 ;
        RECT  2.830 1.030 3.130 1.360 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.420 1.570 8.710 2.540 ;
        RECT  0.260 2.260 0.540 2.880 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  6.260 -0.140 6.420 0.420 ;
        RECT  0.180 -0.140 0.460 0.380 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  6.330 4.260 6.610 4.940 ;
        RECT  2.940 4.260 3.220 4.940 ;
        RECT  1.320 4.270 1.600 4.940 ;
        RECT  0.230 4.280 0.510 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.090 0.740 1.870 0.900 ;
        RECT  0.440 1.080 1.250 1.240 ;
        RECT  1.090 0.740 1.250 1.780 ;
        RECT  1.050 1.080 1.250 1.780 ;
        RECT  1.050 1.550 3.130 1.780 ;
        RECT  1.830 3.020 3.460 3.180 ;
        RECT  3.300 3.020 3.460 3.740 ;
        RECT  1.830 3.020 2.000 3.790 ;
        RECT  1.350 3.510 2.000 3.790 ;
        RECT  1.840 3.020 2.000 4.450 ;
        RECT  1.840 4.290 2.300 4.450 ;
        RECT  3.620 2.700 3.930 2.920 ;
        RECT  3.620 2.700 3.860 3.400 ;
        RECT  3.700 2.700 3.860 4.180 ;
        RECT  3.700 3.910 3.980 4.180 ;
        RECT  0.770 0.300 4.440 0.460 ;
        RECT  4.140 0.300 4.440 0.570 ;
        RECT  0.770 0.300 0.930 0.860 ;
        RECT  0.590 0.580 0.930 0.860 ;
        RECT  0.630 1.780 0.870 2.100 ;
        RECT  4.200 1.890 4.540 2.100 ;
        RECT  0.630 1.940 4.540 2.100 ;
        RECT  4.440 3.020 4.940 3.260 ;
        RECT  2.160 3.450 2.360 4.100 ;
        RECT  2.160 3.940 3.540 4.100 ;
        RECT  3.380 3.940 3.540 4.500 ;
        RECT  4.260 3.980 4.600 4.500 ;
        RECT  4.440 3.020 4.600 4.500 ;
        RECT  3.380 4.340 4.600 4.500 ;
        RECT  4.050 1.070 5.770 1.230 ;
        RECT  4.050 1.070 4.340 1.390 ;
        RECT  5.570 0.620 5.770 1.780 ;
        RECT  5.570 1.620 5.970 1.780 ;
        RECT  5.650 3.020 7.170 3.220 ;
        RECT  6.890 3.020 7.170 3.460 ;
        RECT  5.650 3.020 5.810 4.180 ;
        RECT  5.430 3.880 5.810 4.180 ;
        RECT  3.290 1.550 4.860 1.710 ;
        RECT  3.290 1.550 3.650 1.780 ;
        RECT  4.700 1.550 4.860 2.100 ;
        RECT  4.700 1.940 7.680 2.100 ;
        RECT  6.010 3.940 7.820 4.100 ;
        RECT  4.760 3.420 4.920 4.500 ;
        RECT  6.010 3.940 6.170 4.500 ;
        RECT  4.760 4.340 6.170 4.500 ;
        RECT  6.970 0.640 7.250 1.240 ;
        RECT  6.970 0.960 7.850 1.240 ;
        RECT  6.970 0.640 7.130 1.760 ;
        RECT  6.710 1.500 7.130 1.760 ;
        RECT  5.990 3.500 6.290 3.780 ;
        RECT  5.990 3.620 8.630 3.780 ;
        RECT  8.350 3.340 8.630 4.420 ;
        RECT  8.340 3.620 8.630 4.420 ;
        RECT  4.120 2.700 8.940 2.860 ;
        RECT  5.220 2.700 5.420 3.690 ;
        RECT  4.120 2.700 4.280 3.740 ;
        RECT  4.020 3.340 4.280 3.740 ;
        RECT  7.330 3.020 9.170 3.180 ;
        RECT  7.330 3.020 7.530 3.310 ;
        RECT  8.970 3.020 9.170 3.380 ;
        RECT  5.090 0.300 6.100 0.460 ;
        RECT  6.580 0.300 8.890 0.460 ;
        RECT  5.940 0.300 6.100 0.740 ;
        RECT  8.730 0.300 8.890 0.740 ;
        RECT  6.580 0.300 6.740 0.740 ;
        RECT  5.940 0.580 6.740 0.740 ;
        RECT  8.730 0.580 9.170 0.740 ;
        RECT  3.080 0.620 3.980 0.780 ;
        RECT  5.090 0.300 5.330 0.910 ;
        RECT  3.820 0.750 5.330 0.910 ;
        RECT  7.910 0.620 8.250 0.780 ;
        RECT  8.010 0.620 8.250 1.410 ;
        RECT  8.010 1.250 9.230 1.410 ;
        RECT  8.920 1.250 9.230 1.690 ;
        RECT  8.010 0.620 8.190 1.710 ;
        RECT  7.460 1.490 8.190 1.710 ;
        RECT  9.160 3.570 9.320 4.380 ;
        RECT  8.920 4.220 9.320 4.380 ;
        LAYER VTPH ;
        RECT  2.980 1.210 4.190 3.540 ;
        RECT  6.020 1.160 9.600 3.540 ;
        RECT  0.000 1.260 9.600 3.540 ;
        RECT  0.000 1.260 4.120 3.600 ;
        RECT  0.000 1.260 2.810 3.660 ;
        RECT  8.380 1.140 9.600 3.660 ;
        RECT  7.030 1.160 9.060 3.860 ;
        LAYER VTNH ;
        RECT  2.810 3.600 7.030 4.800 ;
        RECT  4.120 3.540 7.030 4.800 ;
        RECT  0.000 3.660 7.030 4.800 ;
        RECT  9.060 3.660 9.600 4.800 ;
        RECT  0.000 3.860 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  0.000 0.000 8.380 1.160 ;
        RECT  0.000 0.000 6.020 1.210 ;
        RECT  0.000 0.000 2.980 1.260 ;
        RECT  4.190 0.000 6.020 1.260 ;
    END
END SDFEQRM4HM

MACRO SDFEQRM2HM
    CLASS CORE ;
    FOREIGN SDFEQRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.306  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.010 2.700 1.210 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  1.160 1.260 2.830 1.430 ;
        RECT  2.500 0.940 2.830 1.430 ;
        RECT  1.160 1.120 1.440 1.430 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        ANTENNAGATEAREA 0.122  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.441  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.010 3.500 1.210 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.150 0.950 3.520 1.390 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.200 1.130 7.560 1.500 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.060 0.840 6.310 1.350 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.410 2.810 0.700 4.470 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 3.240 2.480 3.690 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.600 0.890 2.320 1.100 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.400 1.690 8.680 2.540 ;
        RECT  2.670 2.260 2.960 2.640 ;
        RECT  0.930 2.260 1.210 3.180 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  6.430 -0.140 6.710 0.320 ;
        RECT  1.840 -0.140 2.120 0.380 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  6.020 4.160 6.180 4.940 ;
        RECT  2.430 4.260 2.710 4.940 ;
        RECT  0.930 4.300 1.210 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.560 0.620 1.310 0.890 ;
        RECT  0.290 0.910 0.740 1.150 ;
        RECT  0.560 0.620 0.740 1.750 ;
        RECT  0.560 1.590 2.810 1.750 ;
        RECT  1.460 2.870 3.030 3.030 ;
        RECT  2.750 2.870 3.030 3.700 ;
        RECT  0.870 3.520 1.620 3.800 ;
        RECT  1.460 2.870 1.620 4.500 ;
        RECT  1.410 3.520 1.620 4.500 ;
        RECT  1.410 4.260 1.690 4.500 ;
        RECT  3.240 2.700 3.520 4.180 ;
        RECT  0.150 1.620 0.400 2.070 ;
        RECT  0.150 1.910 4.230 2.070 ;
        RECT  0.120 0.300 1.680 0.460 ;
        RECT  2.430 0.300 4.350 0.460 ;
        RECT  1.520 0.300 1.680 0.700 ;
        RECT  4.000 0.300 4.350 0.540 ;
        RECT  0.120 0.300 0.400 0.700 ;
        RECT  2.430 0.300 2.590 0.700 ;
        RECT  1.520 0.540 2.590 0.700 ;
        RECT  4.090 3.020 4.860 3.280 ;
        RECT  1.780 3.440 1.940 4.100 ;
        RECT  1.780 3.940 3.030 4.100 ;
        RECT  2.870 3.940 3.030 4.500 ;
        RECT  4.090 3.020 4.340 4.500 ;
        RECT  2.870 4.340 4.340 4.500 ;
        RECT  5.550 0.650 5.900 0.910 ;
        RECT  3.720 1.120 5.710 1.280 ;
        RECT  3.720 1.120 4.020 1.400 ;
        RECT  5.550 0.650 5.710 1.760 ;
        RECT  5.550 1.600 6.030 1.760 ;
        RECT  2.970 1.550 3.290 1.750 ;
        RECT  2.970 1.590 4.790 1.750 ;
        RECT  4.620 1.590 4.790 2.100 ;
        RECT  4.620 1.940 7.540 2.100 ;
        RECT  5.340 3.020 5.620 3.670 ;
        RECT  5.340 3.510 6.820 3.670 ;
        RECT  5.340 3.020 5.520 3.720 ;
        RECT  6.660 3.510 6.820 4.180 ;
        RECT  5.360 3.020 5.520 4.180 ;
        RECT  6.660 3.970 7.820 4.180 ;
        RECT  5.700 3.830 6.500 3.990 ;
        RECT  4.920 4.160 5.200 4.500 ;
        RECT  6.340 3.830 6.500 4.500 ;
        RECT  5.700 3.830 5.860 4.500 ;
        RECT  4.920 4.340 5.860 4.500 ;
        RECT  8.040 3.900 8.200 4.500 ;
        RECT  6.340 4.340 8.200 4.500 ;
        RECT  6.100 3.190 7.140 3.350 ;
        RECT  6.980 3.190 7.140 3.720 ;
        RECT  8.360 3.340 8.640 3.720 ;
        RECT  6.980 3.560 8.640 3.720 ;
        RECT  8.400 3.340 8.640 4.470 ;
        RECT  7.190 0.620 7.980 0.850 ;
        RECT  6.740 0.800 7.440 0.960 ;
        RECT  7.820 0.620 7.980 1.210 ;
        RECT  7.820 0.990 8.730 1.210 ;
        RECT  6.740 0.800 7.020 1.760 ;
        RECT  3.740 2.700 9.010 2.860 ;
        RECT  5.020 2.700 5.180 3.680 ;
        RECT  3.740 2.700 3.900 3.920 ;
        RECT  3.680 3.600 3.900 3.920 ;
        RECT  7.300 3.020 9.240 3.180 ;
        RECT  8.960 3.020 9.240 3.260 ;
        RECT  7.300 3.020 7.560 3.400 ;
        RECT  8.510 0.620 9.270 0.780 ;
        RECT  7.720 1.370 9.270 1.530 ;
        RECT  7.720 1.370 8.030 1.650 ;
        RECT  9.110 0.620 9.270 1.710 ;
        RECT  8.990 1.370 9.270 1.710 ;
        RECT  9.220 3.560 9.500 4.450 ;
        RECT  8.920 4.170 9.500 4.450 ;
        RECT  4.980 0.300 6.220 0.460 ;
        RECT  6.870 0.300 9.500 0.460 ;
        RECT  6.060 0.300 6.220 0.640 ;
        RECT  6.870 0.300 7.030 0.640 ;
        RECT  6.060 0.480 7.030 0.640 ;
        RECT  2.760 0.620 3.850 0.780 ;
        RECT  4.980 0.300 5.140 0.930 ;
        RECT  3.680 0.770 5.140 0.930 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.670 3.660 ;
        RECT  0.000 1.190 9.600 3.540 ;
        RECT  0.000 1.190 3.960 3.610 ;
        RECT  0.000 1.190 1.430 3.660 ;
        RECT  7.930 1.140 9.600 3.660 ;
        RECT  6.650 1.190 9.070 3.860 ;
        LAYER VTNH ;
        RECT  1.430 3.610 6.650 4.800 ;
        RECT  3.960 3.540 6.650 4.800 ;
        RECT  0.000 3.660 6.650 4.800 ;
        RECT  9.070 3.660 9.600 4.800 ;
        RECT  0.000 3.860 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  0.670 0.000 7.930 1.190 ;
    END
END SDFEQRM2HM

MACRO SDFEQRM1HM
    CLASS CORE ;
    FOREIGN SDFEQRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.306  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.010 2.700 1.210 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  1.160 1.260 2.830 1.430 ;
        RECT  2.500 0.940 2.830 1.430 ;
        RECT  1.160 1.120 1.440 1.430 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.545  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.010 3.500 1.210 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.150 0.950 3.520 1.390 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.200 1.130 7.560 1.500 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.060 0.800 6.310 1.350 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.410 2.810 0.700 4.410 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 3.220 2.490 3.570 ;
        END
    END RB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.600 0.890 2.320 1.100 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.400 1.690 8.680 2.540 ;
        RECT  2.670 2.260 2.960 2.640 ;
        RECT  0.930 2.260 1.210 3.030 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  6.430 -0.140 6.710 0.320 ;
        RECT  1.840 -0.140 2.120 0.380 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  6.020 4.160 6.180 4.940 ;
        RECT  2.430 4.260 2.710 4.940 ;
        RECT  0.930 4.300 1.210 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.560 0.620 1.300 0.890 ;
        RECT  0.290 0.910 0.740 1.150 ;
        RECT  0.560 0.620 0.740 1.750 ;
        RECT  0.560 1.590 2.810 1.750 ;
        RECT  1.460 2.870 3.030 3.030 ;
        RECT  2.750 2.870 3.030 3.700 ;
        RECT  0.870 3.520 1.620 3.800 ;
        RECT  1.460 2.870 1.620 4.500 ;
        RECT  1.410 3.520 1.620 4.500 ;
        RECT  1.410 4.260 1.730 4.500 ;
        RECT  3.240 2.700 3.520 4.180 ;
        RECT  0.150 1.620 0.400 2.070 ;
        RECT  0.150 1.910 4.230 2.070 ;
        RECT  0.120 0.300 1.680 0.460 ;
        RECT  2.430 0.300 4.350 0.460 ;
        RECT  1.520 0.300 1.680 0.700 ;
        RECT  4.000 0.300 4.350 0.540 ;
        RECT  0.120 0.300 0.400 0.700 ;
        RECT  2.430 0.300 2.590 0.700 ;
        RECT  1.520 0.540 2.590 0.700 ;
        RECT  4.090 3.020 4.860 3.350 ;
        RECT  1.780 3.440 1.940 4.100 ;
        RECT  1.780 3.940 3.030 4.100 ;
        RECT  2.870 3.940 3.030 4.500 ;
        RECT  4.090 3.020 4.340 4.500 ;
        RECT  2.870 4.340 4.340 4.500 ;
        RECT  5.550 0.650 5.900 0.910 ;
        RECT  3.720 1.120 5.710 1.280 ;
        RECT  3.720 1.120 4.020 1.400 ;
        RECT  5.550 0.650 5.710 1.760 ;
        RECT  5.550 1.600 6.030 1.760 ;
        RECT  2.970 1.550 3.290 1.750 ;
        RECT  2.970 1.590 4.790 1.750 ;
        RECT  4.620 1.590 4.790 2.100 ;
        RECT  4.620 1.940 7.540 2.100 ;
        RECT  5.340 3.020 5.620 3.670 ;
        RECT  5.340 3.510 6.820 3.670 ;
        RECT  5.340 3.020 5.520 3.720 ;
        RECT  6.660 3.510 6.820 4.180 ;
        RECT  5.360 3.020 5.520 4.180 ;
        RECT  6.660 3.970 7.820 4.180 ;
        RECT  5.700 3.830 6.500 3.990 ;
        RECT  4.920 4.160 5.200 4.500 ;
        RECT  6.340 3.830 6.500 4.500 ;
        RECT  5.700 3.830 5.860 4.500 ;
        RECT  4.920 4.340 5.860 4.500 ;
        RECT  8.040 3.900 8.200 4.500 ;
        RECT  6.340 4.340 8.200 4.500 ;
        RECT  6.100 3.190 7.140 3.350 ;
        RECT  6.980 3.190 7.140 3.720 ;
        RECT  8.360 3.340 8.640 3.720 ;
        RECT  6.980 3.560 8.640 3.720 ;
        RECT  8.400 3.340 8.640 4.470 ;
        RECT  7.190 0.620 7.980 0.850 ;
        RECT  6.740 0.800 7.440 0.960 ;
        RECT  7.820 0.620 7.980 1.210 ;
        RECT  7.820 0.990 8.730 1.210 ;
        RECT  6.740 0.800 7.020 1.760 ;
        RECT  3.740 2.700 9.010 2.860 ;
        RECT  5.020 2.700 5.180 3.680 ;
        RECT  3.740 2.700 3.900 3.920 ;
        RECT  3.680 3.600 3.900 3.920 ;
        RECT  7.300 3.020 9.240 3.180 ;
        RECT  8.960 3.020 9.240 3.260 ;
        RECT  7.300 3.020 7.560 3.400 ;
        RECT  8.510 0.620 9.270 0.780 ;
        RECT  7.720 1.370 9.270 1.530 ;
        RECT  7.720 1.370 8.030 1.650 ;
        RECT  9.110 0.620 9.270 1.710 ;
        RECT  8.990 1.370 9.270 1.710 ;
        RECT  9.220 3.560 9.500 4.450 ;
        RECT  8.920 4.170 9.500 4.450 ;
        RECT  5.070 0.300 6.220 0.460 ;
        RECT  6.870 0.300 9.500 0.460 ;
        RECT  6.060 0.300 6.220 0.640 ;
        RECT  6.870 0.300 7.030 0.640 ;
        RECT  6.060 0.480 7.030 0.640 ;
        RECT  2.760 0.620 3.850 0.780 ;
        RECT  5.070 0.300 5.230 0.930 ;
        RECT  3.680 0.770 5.230 0.930 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.670 3.660 ;
        RECT  0.000 1.190 9.600 3.540 ;
        RECT  0.000 1.190 3.960 3.610 ;
        RECT  0.000 1.190 1.430 3.660 ;
        RECT  7.930 1.140 9.600 3.660 ;
        RECT  6.650 1.190 9.070 3.860 ;
        LAYER VTNH ;
        RECT  1.430 3.610 6.650 4.800 ;
        RECT  3.960 3.540 6.650 4.800 ;
        RECT  0.000 3.660 6.650 4.800 ;
        RECT  9.070 3.660 9.600 4.800 ;
        RECT  0.000 3.860 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  0.670 0.000 7.930 1.190 ;
    END
END SDFEQRM1HM

MACRO SDFEQM8HM
    CLASS CORE ;
    FOREIGN SDFEQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.539  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.250 3.420 5.450 3.620 ;
        LAYER ME2 ;
        RECT  5.250 3.240 5.500 3.960 ;
        LAYER ME1 ;
        RECT  5.130 3.340 5.450 3.750 ;
        RECT  5.130 3.340 5.400 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.210 1.610 3.600 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.155  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.530 0.710 4.250 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.236  LAYER ME1  ;
        ANTENNADIFFAREA 1.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.710 0.840 9.160 1.160 ;
        RECT  8.710 0.330 8.990 2.100 ;
        RECT  8.640 0.330 8.990 0.830 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.640 1.010 1.280 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.190 1.490 9.470 3.320 ;
        RECT  8.150 1.500 8.430 3.320 ;
        RECT  7.170 2.260 7.370 3.000 ;
        RECT  6.400 2.120 6.680 2.540 ;
        RECT  5.320 1.700 5.600 2.540 ;
        RECT  3.030 1.770 3.310 2.540 ;
        RECT  2.970 2.260 3.270 3.040 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.040 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.190 -0.140 9.470 0.620 ;
        RECT  8.150 -0.140 8.430 0.610 ;
        RECT  6.120 -0.140 6.400 0.500 ;
        RECT  4.940 -0.140 5.210 0.560 ;
        RECT  2.500 -0.140 2.780 0.320 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  9.200 4.050 9.470 4.940 ;
        RECT  8.190 4.020 8.430 4.940 ;
        RECT  7.090 4.270 7.370 4.940 ;
        RECT  4.770 4.480 5.050 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.200 1.030 3.370 ;
        RECT  0.870 3.200 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.040 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.640 1.130 2.560 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.640 1.130 1.800 1.820 ;
        RECT  0.100 1.660 1.800 1.820 ;
        RECT  1.070 0.300 2.240 0.460 ;
        RECT  2.070 0.300 2.240 0.640 ;
        RECT  3.100 0.320 3.380 0.640 ;
        RECT  2.070 0.480 3.380 0.640 ;
        RECT  1.070 0.300 1.310 0.830 ;
        RECT  1.570 0.620 1.850 0.960 ;
        RECT  3.580 0.340 3.860 0.960 ;
        RECT  1.570 0.800 3.860 0.960 ;
        RECT  3.610 2.700 3.970 2.960 ;
        RECT  3.610 2.700 3.790 4.160 ;
        RECT  3.350 3.940 3.790 4.160 ;
        RECT  2.710 1.410 4.010 1.610 ;
        RECT  2.070 1.600 2.870 1.770 ;
        RECT  4.770 3.020 5.920 3.180 ;
        RECT  5.610 3.020 5.920 3.720 ;
        RECT  4.770 3.020 4.930 3.660 ;
        RECT  4.590 3.440 4.930 3.660 ;
        RECT  5.610 3.430 6.000 3.720 ;
        RECT  5.610 3.020 5.850 4.150 ;
        RECT  5.560 3.900 5.850 4.150 ;
        RECT  4.090 0.340 4.420 0.670 ;
        RECT  4.240 0.340 4.420 1.650 ;
        RECT  4.240 1.040 6.200 1.200 ;
        RECT  4.240 1.040 4.520 1.650 ;
        RECT  4.190 2.700 6.580 2.860 ;
        RECT  4.190 2.700 4.350 3.360 ;
        RECT  3.950 3.120 4.230 4.150 ;
        RECT  6.360 1.040 7.340 1.320 ;
        RECT  6.360 1.040 6.520 1.520 ;
        RECT  4.810 1.360 6.520 1.520 ;
        RECT  4.810 1.360 4.970 2.040 ;
        RECT  3.480 1.810 4.970 2.040 ;
        RECT  6.130 3.080 6.410 3.300 ;
        RECT  6.160 3.160 7.430 3.320 ;
        RECT  7.270 3.160 7.430 3.750 ;
        RECT  7.270 3.500 7.550 3.750 ;
        RECT  6.160 3.160 6.440 4.180 ;
        RECT  6.100 3.900 6.440 4.180 ;
        RECT  5.600 0.460 5.880 0.880 ;
        RECT  6.640 0.340 6.920 0.880 ;
        RECT  4.720 0.720 7.670 0.880 ;
        RECT  7.510 0.720 7.670 1.640 ;
        RECT  7.140 1.480 7.670 1.640 ;
        RECT  5.800 1.680 7.320 1.840 ;
        RECT  7.140 1.480 7.320 1.860 ;
        RECT  6.970 1.660 7.320 1.860 ;
        RECT  7.690 2.700 7.890 3.030 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  6.760 3.510 7.070 4.070 ;
        RECT  6.760 3.910 7.890 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.450 4.160 5.370 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.210 4.160 5.370 4.500 ;
        RECT  7.710 2.700 7.890 4.490 ;
        RECT  7.630 3.910 7.890 4.490 ;
        RECT  4.450 4.160 4.610 4.500 ;
        RECT  3.030 4.340 4.610 4.500 ;
        RECT  6.760 3.510 6.920 4.500 ;
        RECT  5.210 4.340 6.920 4.500 ;
        RECT  7.160 0.340 7.990 0.500 ;
        RECT  7.830 1.030 8.490 1.250 ;
        RECT  7.830 0.340 7.990 1.960 ;
        RECT  7.480 1.800 7.990 1.960 ;
        RECT  8.670 2.740 8.950 4.470 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 3.540 ;
        RECT  3.460 1.070 7.980 3.600 ;
        RECT  2.860 1.140 9.600 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.330 1.140 9.600 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.330 4.800 ;
        RECT  0.000 3.660 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.070 ;
        RECT  0.000 0.000 3.460 1.140 ;
        RECT  7.980 0.000 9.600 1.140 ;
    END
END SDFEQM8HM

MACRO SDFEQM4HM
    CLASS CORE ;
    FOREIGN SDFEQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.635  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.280 3.420 5.480 3.620 ;
        LAYER ME2 ;
        RECT  5.280 3.240 5.530 3.960 ;
        LAYER ME1 ;
        RECT  5.160 3.340 5.480 3.750 ;
        RECT  5.160 3.340 5.430 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.220 1.610 3.600 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.540 0.710 4.310 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.158  LAYER ME1  ;
        ANTENNADIFFAREA 0.933  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.800 0.840 9.100 1.210 ;
        RECT  8.800 0.330 9.080 2.100 ;
        RECT  8.730 0.330 9.080 0.830 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.010 1.320 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.240 1.500 8.520 3.330 ;
        RECT  7.200 2.260 7.400 3.000 ;
        RECT  5.430 1.680 5.710 2.540 ;
        RECT  3.110 1.770 3.390 2.540 ;
        RECT  2.970 2.260 3.270 3.050 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.050 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.240 -0.140 8.520 0.610 ;
        RECT  5.190 -0.140 5.460 0.560 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  0.000 4.660 9.200 4.940 ;
        RECT  8.280 4.020 8.520 4.940 ;
        RECT  7.160 4.300 7.440 4.940 ;
        RECT  4.800 4.480 5.080 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.210 1.030 3.380 ;
        RECT  0.870 3.210 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.050 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.720 1.130 2.640 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.720 1.130 1.880 1.820 ;
        RECT  0.100 1.660 1.880 1.820 ;
        RECT  1.010 0.300 2.320 0.460 ;
        RECT  2.150 0.300 2.320 0.640 ;
        RECT  3.180 0.320 3.460 0.640 ;
        RECT  2.150 0.480 3.460 0.640 ;
        RECT  1.010 0.300 1.290 0.830 ;
        RECT  1.650 0.620 1.930 0.960 ;
        RECT  3.690 0.340 3.970 0.960 ;
        RECT  1.650 0.800 3.970 0.960 ;
        RECT  3.640 2.700 4.000 2.960 ;
        RECT  3.640 2.700 3.820 4.160 ;
        RECT  3.350 3.940 3.820 4.160 ;
        RECT  2.790 1.410 4.120 1.610 ;
        RECT  2.150 1.600 2.950 1.770 ;
        RECT  4.200 0.340 4.670 0.670 ;
        RECT  4.350 0.340 4.670 1.200 ;
        RECT  4.350 1.040 5.880 1.200 ;
        RECT  4.350 0.340 4.590 1.650 ;
        RECT  4.800 3.020 5.950 3.180 ;
        RECT  5.640 3.020 5.950 3.720 ;
        RECT  4.800 3.020 4.960 3.660 ;
        RECT  4.620 3.440 4.960 3.660 ;
        RECT  5.640 3.430 6.030 3.720 ;
        RECT  5.640 3.020 5.880 4.150 ;
        RECT  5.590 3.900 5.880 4.150 ;
        RECT  4.220 2.700 6.700 2.860 ;
        RECT  4.220 2.700 4.380 3.360 ;
        RECT  3.980 3.120 4.260 4.150 ;
        RECT  6.040 1.040 7.010 1.320 ;
        RECT  6.040 1.040 6.200 1.520 ;
        RECT  4.920 1.360 6.200 1.520 ;
        RECT  4.920 1.360 5.080 2.040 ;
        RECT  3.590 1.810 5.080 2.040 ;
        RECT  5.710 0.460 5.990 0.880 ;
        RECT  6.310 0.340 6.590 0.880 ;
        RECT  4.830 0.720 7.340 0.880 ;
        RECT  7.180 0.720 7.340 1.640 ;
        RECT  6.810 1.480 7.340 1.640 ;
        RECT  5.910 1.680 6.990 1.840 ;
        RECT  6.810 1.480 6.990 1.860 ;
        RECT  6.640 1.660 6.990 1.860 ;
        RECT  6.160 3.080 6.440 3.300 ;
        RECT  6.190 3.160 7.460 3.320 ;
        RECT  7.300 3.160 7.460 3.750 ;
        RECT  7.300 3.500 7.620 3.750 ;
        RECT  6.190 3.160 6.470 4.180 ;
        RECT  6.130 3.900 6.470 4.180 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  6.790 3.510 7.140 4.070 ;
        RECT  6.790 3.910 8.040 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.480 4.160 5.400 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.240 4.160 5.400 4.500 ;
        RECT  7.800 2.700 8.040 4.490 ;
        RECT  7.760 3.910 8.040 4.490 ;
        RECT  4.480 4.160 4.640 4.500 ;
        RECT  3.030 4.340 4.640 4.500 ;
        RECT  6.790 3.510 6.950 4.500 ;
        RECT  5.240 4.340 6.950 4.500 ;
        RECT  6.910 0.340 7.720 0.500 ;
        RECT  7.560 1.030 8.580 1.250 ;
        RECT  7.560 0.340 7.720 1.960 ;
        RECT  7.150 1.800 7.720 1.960 ;
        RECT  8.760 2.740 9.040 4.470 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.200 3.540 ;
        RECT  3.570 1.070 7.650 3.600 ;
        RECT  2.860 1.140 9.200 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.360 1.140 9.200 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.360 4.800 ;
        RECT  0.000 3.660 9.200 4.800 ;
        RECT  0.000 0.000 9.200 1.070 ;
        RECT  0.000 0.000 3.570 1.140 ;
        RECT  7.650 0.000 9.200 1.140 ;
    END
END SDFEQM4HM

MACRO SDFEQM2HM
    CLASS CORE ;
    FOREIGN SDFEQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.240 3.340 5.660 3.750 ;
        RECT  5.240 3.340 5.610 3.960 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.220 1.610 3.600 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.540 0.710 4.310 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.380 0.840 8.700 1.210 ;
        RECT  8.380 0.330 8.620 2.100 ;
        RECT  8.310 0.330 8.620 0.830 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.010 1.280 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.820 1.500 8.100 2.540 ;
        RECT  7.380 2.260 7.580 3.000 ;
        RECT  5.430 1.680 5.710 2.540 ;
        RECT  3.110 1.770 3.390 2.540 ;
        RECT  2.970 2.260 3.270 3.050 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.050 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.820 -0.140 8.100 0.610 ;
        RECT  5.190 -0.140 5.460 0.560 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  0.000 4.660 8.800 4.940 ;
        RECT  7.340 4.300 7.620 4.940 ;
        RECT  4.800 4.480 5.080 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.210 1.030 3.380 ;
        RECT  0.870 3.210 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.050 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.720 1.130 2.640 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.720 1.130 1.880 1.820 ;
        RECT  0.100 1.660 1.880 1.820 ;
        RECT  1.010 0.300 2.320 0.460 ;
        RECT  2.150 0.300 2.320 0.640 ;
        RECT  3.180 0.320 3.460 0.640 ;
        RECT  2.150 0.480 3.460 0.640 ;
        RECT  1.010 0.300 1.290 0.820 ;
        RECT  1.650 0.620 1.930 0.960 ;
        RECT  3.690 0.340 3.970 0.960 ;
        RECT  1.650 0.800 3.970 0.960 ;
        RECT  3.640 2.700 4.000 2.960 ;
        RECT  3.640 2.700 3.820 4.160 ;
        RECT  3.350 3.940 3.820 4.160 ;
        RECT  2.790 1.410 4.120 1.610 ;
        RECT  2.150 1.600 2.950 1.770 ;
        RECT  4.200 0.340 4.670 0.670 ;
        RECT  4.350 0.340 4.670 1.200 ;
        RECT  4.350 1.040 5.880 1.200 ;
        RECT  4.350 0.340 4.590 1.650 ;
        RECT  4.800 3.020 6.130 3.180 ;
        RECT  5.820 3.020 6.130 3.720 ;
        RECT  4.800 3.020 4.960 3.660 ;
        RECT  4.620 3.440 4.960 3.660 ;
        RECT  5.820 3.430 6.210 3.720 ;
        RECT  5.820 3.020 6.060 4.150 ;
        RECT  5.770 3.900 6.060 4.150 ;
        RECT  4.220 2.700 6.880 2.860 ;
        RECT  4.220 2.700 4.380 3.360 ;
        RECT  3.980 3.120 4.260 4.150 ;
        RECT  6.040 1.040 7.010 1.320 ;
        RECT  6.040 1.040 6.200 1.520 ;
        RECT  4.920 1.360 6.200 1.520 ;
        RECT  4.920 1.360 5.080 2.040 ;
        RECT  3.590 1.810 5.080 2.040 ;
        RECT  5.710 0.460 5.990 0.880 ;
        RECT  6.310 0.340 6.590 0.880 ;
        RECT  4.910 0.720 7.340 0.880 ;
        RECT  7.180 0.720 7.340 1.640 ;
        RECT  6.810 1.480 7.340 1.640 ;
        RECT  5.910 1.680 6.990 1.840 ;
        RECT  6.810 1.480 6.990 1.860 ;
        RECT  6.640 1.660 6.990 1.860 ;
        RECT  6.340 3.080 6.620 3.300 ;
        RECT  6.370 3.160 7.640 3.320 ;
        RECT  7.480 3.160 7.640 3.750 ;
        RECT  7.480 3.500 7.800 3.750 ;
        RECT  6.370 3.160 6.650 4.180 ;
        RECT  6.310 3.900 6.650 4.180 ;
        RECT  6.910 0.340 7.660 0.500 ;
        RECT  7.500 1.030 8.160 1.250 ;
        RECT  7.500 0.340 7.660 1.960 ;
        RECT  7.150 1.800 7.660 1.960 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  6.970 3.510 7.320 4.070 ;
        RECT  6.970 3.910 8.220 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.480 4.160 5.580 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.420 4.160 5.580 4.500 ;
        RECT  7.980 2.700 8.220 4.490 ;
        RECT  7.940 3.910 8.220 4.490 ;
        RECT  4.480 4.160 4.640 4.500 ;
        RECT  3.030 4.340 4.640 4.500 ;
        RECT  6.970 3.510 7.130 4.500 ;
        RECT  5.420 4.340 7.130 4.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 3.540 ;
        RECT  3.570 1.070 7.590 3.600 ;
        RECT  2.860 1.140 8.800 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.540 1.140 8.800 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.540 4.800 ;
        RECT  0.000 3.660 8.800 4.800 ;
        RECT  0.000 0.000 8.800 1.070 ;
        RECT  0.000 0.000 3.570 1.140 ;
        RECT  7.590 0.000 8.800 1.140 ;
    END
END SDFEQM2HM

MACRO SDFEQM1HM
    CLASS CORE ;
    FOREIGN SDFEQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.240 3.340 5.660 3.750 ;
        RECT  5.240 3.340 5.610 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.220 1.610 3.600 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.150  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.540 0.710 4.310 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.380 0.840 8.700 1.210 ;
        RECT  8.380 0.300 8.620 2.100 ;
        RECT  8.310 0.300 8.620 0.830 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.010 1.280 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.820 1.760 8.100 2.540 ;
        RECT  7.380 2.260 7.580 3.000 ;
        RECT  5.430 1.680 5.710 2.540 ;
        RECT  3.110 1.770 3.390 2.540 ;
        RECT  2.970 2.260 3.270 3.050 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.050 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.820 -0.140 8.100 0.610 ;
        RECT  5.190 -0.140 5.460 0.560 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  0.000 4.660 8.800 4.940 ;
        RECT  7.340 4.300 7.620 4.940 ;
        RECT  4.800 4.480 5.080 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.210 1.030 3.380 ;
        RECT  0.870 3.210 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.050 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.720 1.130 2.640 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.720 1.130 1.880 1.820 ;
        RECT  0.100 1.660 1.880 1.820 ;
        RECT  1.010 0.300 2.320 0.460 ;
        RECT  2.150 0.300 2.320 0.640 ;
        RECT  3.180 0.320 3.460 0.640 ;
        RECT  2.150 0.480 3.460 0.640 ;
        RECT  1.010 0.300 1.290 0.830 ;
        RECT  1.650 0.620 1.930 0.960 ;
        RECT  3.690 0.340 3.970 0.960 ;
        RECT  1.650 0.800 3.970 0.960 ;
        RECT  3.640 2.700 4.000 2.960 ;
        RECT  3.640 2.700 3.820 4.160 ;
        RECT  3.350 3.940 3.820 4.160 ;
        RECT  2.790 1.410 4.120 1.610 ;
        RECT  2.150 1.600 2.950 1.770 ;
        RECT  4.200 0.340 4.670 0.670 ;
        RECT  4.350 0.340 4.670 1.200 ;
        RECT  4.350 1.040 5.880 1.200 ;
        RECT  4.350 0.340 4.590 1.650 ;
        RECT  4.800 3.020 6.130 3.180 ;
        RECT  5.820 3.020 6.130 3.720 ;
        RECT  4.800 3.020 4.960 3.660 ;
        RECT  4.620 3.440 4.960 3.660 ;
        RECT  5.820 3.430 6.210 3.720 ;
        RECT  5.820 3.020 6.060 4.150 ;
        RECT  5.770 3.900 6.060 4.150 ;
        RECT  4.220 2.700 6.880 2.860 ;
        RECT  4.220 2.700 4.380 3.360 ;
        RECT  3.980 3.120 4.260 4.150 ;
        RECT  6.040 1.040 7.010 1.320 ;
        RECT  6.040 1.040 6.200 1.520 ;
        RECT  4.920 1.360 6.200 1.520 ;
        RECT  4.920 1.360 5.080 2.040 ;
        RECT  3.590 1.810 5.080 2.040 ;
        RECT  5.710 0.460 5.990 0.880 ;
        RECT  6.310 0.340 6.590 0.880 ;
        RECT  4.830 0.720 7.340 0.880 ;
        RECT  7.180 0.720 7.340 1.640 ;
        RECT  6.810 1.480 7.340 1.640 ;
        RECT  5.910 1.680 6.990 1.840 ;
        RECT  6.810 1.480 6.990 1.860 ;
        RECT  6.640 1.660 6.990 1.860 ;
        RECT  6.340 3.080 6.620 3.300 ;
        RECT  6.370 3.160 7.640 3.320 ;
        RECT  7.480 3.160 7.640 3.750 ;
        RECT  7.480 3.500 7.800 3.750 ;
        RECT  6.370 3.160 6.650 4.180 ;
        RECT  6.310 3.900 6.650 4.180 ;
        RECT  6.910 0.340 7.660 0.500 ;
        RECT  7.500 1.030 8.160 1.250 ;
        RECT  7.500 0.340 7.660 1.960 ;
        RECT  7.150 1.800 7.660 1.960 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  6.970 3.510 7.320 4.070 ;
        RECT  6.970 3.910 8.220 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.480 4.160 5.580 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.420 4.160 5.580 4.500 ;
        RECT  7.980 2.700 8.220 4.490 ;
        RECT  7.940 3.910 8.220 4.490 ;
        RECT  4.480 4.160 4.640 4.500 ;
        RECT  3.030 4.340 4.640 4.500 ;
        RECT  6.970 3.510 7.130 4.500 ;
        RECT  5.420 4.340 7.130 4.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 3.540 ;
        RECT  3.570 1.070 7.590 3.600 ;
        RECT  2.860 1.140 8.800 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.540 1.140 8.800 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.540 4.800 ;
        RECT  0.000 3.660 8.800 4.800 ;
        RECT  0.000 0.000 8.800 1.070 ;
        RECT  0.000 0.000 3.570 1.140 ;
        RECT  7.590 0.000 8.800 1.140 ;
    END
END SDFEQM1HM

MACRO SDFEM8HM
    CLASS CORE ;
    FOREIGN SDFEM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.539  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.250 3.420 5.450 3.620 ;
        LAYER ME2 ;
        RECT  5.250 3.240 5.500 3.960 ;
        LAYER ME1 ;
        RECT  5.130 3.340 5.450 3.750 ;
        RECT  5.130 3.340 5.400 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.210 1.610 3.600 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.155  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.530 0.710 4.250 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.750 0.480 10.030 2.100 ;
        RECT  8.710 0.900 10.030 1.210 ;
        RECT  9.680 0.480 10.030 1.210 ;
        RECT  8.710 0.480 8.990 2.100 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.710 2.740 9.990 4.470 ;
        RECT  8.670 3.530 9.990 3.900 ;
        RECT  8.670 2.740 8.950 4.470 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.000 1.290 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  10.230 1.490 10.510 3.330 ;
        RECT  9.190 1.490 9.470 3.330 ;
        RECT  8.150 1.500 8.430 3.330 ;
        RECT  7.170 2.260 7.370 3.000 ;
        RECT  6.400 2.120 6.680 2.540 ;
        RECT  5.320 1.700 5.600 2.540 ;
        RECT  3.030 1.770 3.310 2.540 ;
        RECT  2.970 2.260 3.270 3.040 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.040 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  10.230 -0.140 10.510 0.710 ;
        RECT  9.190 -0.140 9.470 0.710 ;
        RECT  8.150 -0.140 8.430 0.610 ;
        RECT  6.120 -0.140 6.400 0.500 ;
        RECT  4.940 -0.140 5.210 0.560 ;
        RECT  2.500 -0.140 2.780 0.320 ;
        RECT  0.000 4.660 10.800 4.940 ;
        RECT  10.240 4.050 10.510 4.940 ;
        RECT  9.190 4.120 9.470 4.940 ;
        RECT  8.190 4.020 8.430 4.940 ;
        RECT  7.090 4.270 7.370 4.940 ;
        RECT  4.770 4.480 5.050 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.200 1.030 3.370 ;
        RECT  0.870 3.200 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.040 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.640 1.130 2.560 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.640 1.130 1.800 1.820 ;
        RECT  0.100 1.660 1.800 1.820 ;
        RECT  1.070 0.300 2.240 0.460 ;
        RECT  2.070 0.300 2.240 0.640 ;
        RECT  3.100 0.320 3.380 0.640 ;
        RECT  2.070 0.480 3.380 0.640 ;
        RECT  1.070 0.300 1.310 0.830 ;
        RECT  1.570 0.620 1.850 0.960 ;
        RECT  3.580 0.340 3.860 0.960 ;
        RECT  1.570 0.800 3.860 0.960 ;
        RECT  3.610 2.700 3.970 2.960 ;
        RECT  3.610 2.700 3.790 4.160 ;
        RECT  3.350 3.940 3.790 4.160 ;
        RECT  2.710 1.410 4.010 1.610 ;
        RECT  2.070 1.600 2.870 1.770 ;
        RECT  4.770 3.020 5.920 3.180 ;
        RECT  5.610 3.020 5.920 3.720 ;
        RECT  4.770 3.020 4.930 3.660 ;
        RECT  4.590 3.440 4.930 3.660 ;
        RECT  5.610 3.430 6.000 3.720 ;
        RECT  5.610 3.020 5.850 4.150 ;
        RECT  5.560 3.900 5.850 4.150 ;
        RECT  4.090 0.340 4.560 0.670 ;
        RECT  4.240 0.340 4.560 1.200 ;
        RECT  4.240 1.040 6.200 1.200 ;
        RECT  4.240 0.340 4.480 1.650 ;
        RECT  4.190 2.700 6.580 2.860 ;
        RECT  4.190 2.700 4.350 3.360 ;
        RECT  3.950 3.120 4.230 4.150 ;
        RECT  6.360 1.040 7.340 1.320 ;
        RECT  6.360 1.040 6.520 1.520 ;
        RECT  4.810 1.360 6.520 1.520 ;
        RECT  4.810 1.360 4.970 2.040 ;
        RECT  3.480 1.810 4.970 2.040 ;
        RECT  6.130 3.080 6.410 3.300 ;
        RECT  6.160 3.160 7.390 3.320 ;
        RECT  7.230 3.160 7.390 3.750 ;
        RECT  7.230 3.500 7.570 3.750 ;
        RECT  6.160 3.160 6.440 4.180 ;
        RECT  6.100 3.900 6.440 4.180 ;
        RECT  5.600 0.460 5.880 0.880 ;
        RECT  6.640 0.340 6.920 0.880 ;
        RECT  4.720 0.720 7.670 0.880 ;
        RECT  7.510 0.720 7.670 1.660 ;
        RECT  7.140 1.500 7.670 1.660 ;
        RECT  5.800 1.680 7.320 1.840 ;
        RECT  7.140 1.500 7.320 1.880 ;
        RECT  6.970 1.680 7.320 1.880 ;
        RECT  7.690 2.700 7.890 3.070 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  7.730 3.510 8.430 3.790 ;
        RECT  6.760 3.510 7.070 4.070 ;
        RECT  6.760 3.910 7.890 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.450 4.160 5.370 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.210 4.160 5.370 4.500 ;
        RECT  7.730 2.700 7.890 4.490 ;
        RECT  7.630 3.910 7.890 4.490 ;
        RECT  4.450 4.160 4.610 4.500 ;
        RECT  3.030 4.340 4.610 4.500 ;
        RECT  6.760 3.510 6.920 4.500 ;
        RECT  5.210 4.340 6.920 4.500 ;
        RECT  7.160 0.340 7.990 0.500 ;
        RECT  7.830 1.030 8.490 1.250 ;
        RECT  7.830 0.340 7.990 1.980 ;
        RECT  7.480 1.820 7.990 1.980 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.800 3.540 ;
        RECT  3.460 1.070 7.950 3.600 ;
        RECT  2.860 1.140 10.800 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.330 1.140 10.800 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.330 4.800 ;
        RECT  0.000 3.660 10.800 4.800 ;
        RECT  0.000 0.000 10.800 1.070 ;
        RECT  0.000 0.000 3.460 1.140 ;
        RECT  7.950 0.000 10.800 1.140 ;
    END
END SDFEM8HM

MACRO SDFEM4HM
    CLASS CORE ;
    FOREIGN SDFEM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.635  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.250 3.420 5.450 3.620 ;
        LAYER ME2 ;
        RECT  5.250 3.240 5.500 3.960 ;
        LAYER ME1 ;
        RECT  5.130 3.340 5.450 3.750 ;
        RECT  5.130 3.340 5.400 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.220 1.610 3.660 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.540 0.710 4.310 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.730 0.840 9.500 1.210 ;
        RECT  8.730 0.330 9.010 2.100 ;
        RECT  8.660 0.330 9.010 0.830 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.690 3.530 9.500 3.960 ;
        RECT  8.690 2.740 8.970 4.470 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.000 1.280 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.210 1.490 9.490 3.330 ;
        RECT  8.170 1.500 8.450 3.330 ;
        RECT  7.210 2.260 7.410 3.000 ;
        RECT  5.320 1.680 5.600 2.540 ;
        RECT  3.030 1.770 3.310 2.540 ;
        RECT  2.970 2.260 3.270 3.050 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.050 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.210 -0.140 9.490 0.650 ;
        RECT  8.170 -0.140 8.450 0.610 ;
        RECT  5.080 -0.140 5.350 0.560 ;
        RECT  2.500 -0.140 2.780 0.320 ;
        RECT  0.000 4.660 9.600 4.940 ;
        RECT  9.210 4.120 9.490 4.940 ;
        RECT  8.210 4.020 8.450 4.940 ;
        RECT  7.130 4.300 7.410 4.940 ;
        RECT  4.770 4.480 5.050 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.210 1.030 3.380 ;
        RECT  0.870 3.210 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.050 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.640 1.130 2.560 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.640 1.130 1.800 1.820 ;
        RECT  0.100 1.660 1.800 1.820 ;
        RECT  1.070 0.300 2.240 0.460 ;
        RECT  2.070 0.300 2.240 0.640 ;
        RECT  3.100 0.320 3.380 0.640 ;
        RECT  2.070 0.480 3.380 0.640 ;
        RECT  1.070 0.300 1.310 0.830 ;
        RECT  1.570 0.620 1.850 0.960 ;
        RECT  3.580 0.340 3.860 0.960 ;
        RECT  1.570 0.800 3.860 0.960 ;
        RECT  3.610 2.700 3.970 2.960 ;
        RECT  3.610 2.700 3.790 4.160 ;
        RECT  3.350 3.940 3.790 4.160 ;
        RECT  2.710 1.410 4.010 1.610 ;
        RECT  2.070 1.600 2.870 1.770 ;
        RECT  4.090 0.340 4.560 0.670 ;
        RECT  4.240 0.340 4.560 1.200 ;
        RECT  4.240 1.040 5.770 1.200 ;
        RECT  4.240 0.340 4.480 1.650 ;
        RECT  4.770 3.020 5.920 3.180 ;
        RECT  5.610 3.020 5.920 3.720 ;
        RECT  4.770 3.020 4.930 3.660 ;
        RECT  4.590 3.440 4.930 3.660 ;
        RECT  5.610 3.430 6.000 3.720 ;
        RECT  5.610 3.020 5.850 4.150 ;
        RECT  5.560 3.900 5.850 4.150 ;
        RECT  4.190 2.700 6.670 2.860 ;
        RECT  4.190 2.700 4.350 3.360 ;
        RECT  3.950 3.120 4.230 4.150 ;
        RECT  5.930 1.040 6.900 1.320 ;
        RECT  5.930 1.040 6.090 1.520 ;
        RECT  4.810 1.360 6.090 1.520 ;
        RECT  4.810 1.360 4.970 2.040 ;
        RECT  3.480 1.810 4.970 2.040 ;
        RECT  5.600 0.460 5.880 0.880 ;
        RECT  6.200 0.340 6.480 0.880 ;
        RECT  4.720 0.720 7.230 0.880 ;
        RECT  7.070 0.720 7.230 1.640 ;
        RECT  6.700 1.480 7.230 1.640 ;
        RECT  5.800 1.680 6.880 1.840 ;
        RECT  6.700 1.480 6.880 1.860 ;
        RECT  6.530 1.660 6.880 1.860 ;
        RECT  6.130 3.080 6.410 3.300 ;
        RECT  6.160 3.160 7.430 3.320 ;
        RECT  7.270 3.160 7.430 3.750 ;
        RECT  7.270 3.500 7.610 3.750 ;
        RECT  6.160 3.160 6.440 4.180 ;
        RECT  6.100 3.900 6.440 4.180 ;
        RECT  7.730 2.700 7.930 3.390 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  7.770 3.510 8.450 3.790 ;
        RECT  6.760 3.510 7.110 4.070 ;
        RECT  6.760 3.910 7.930 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.450 4.160 5.370 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.210 4.160 5.370 4.500 ;
        RECT  7.770 2.700 7.930 4.490 ;
        RECT  7.650 3.910 7.930 4.490 ;
        RECT  4.450 4.160 4.610 4.500 ;
        RECT  3.030 4.340 4.610 4.500 ;
        RECT  6.760 3.510 6.920 4.500 ;
        RECT  5.210 4.340 6.920 4.500 ;
        RECT  6.800 0.340 7.550 0.500 ;
        RECT  7.390 1.030 8.510 1.250 ;
        RECT  7.390 0.340 7.550 1.960 ;
        RECT  7.040 1.800 7.550 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 3.540 ;
        RECT  3.460 1.070 7.540 3.600 ;
        RECT  2.860 1.140 9.600 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.330 1.140 9.600 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.330 4.800 ;
        RECT  0.000 3.660 9.600 4.800 ;
        RECT  0.000 0.000 9.600 1.070 ;
        RECT  0.000 0.000 3.460 1.140 ;
        RECT  7.540 0.000 9.600 1.140 ;
    END
END SDFEM4HM

MACRO SDFEM2HM
    CLASS CORE ;
    FOREIGN SDFEM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.224  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.250 3.420 5.450 3.620 ;
        LAYER ME2 ;
        RECT  5.250 3.240 5.500 3.960 ;
        LAYER ME1 ;
        RECT  5.130 3.340 5.450 3.750 ;
        RECT  4.600 3.830 5.400 4.000 ;
        RECT  5.130 3.340 5.400 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.220 1.610 3.640 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.540 0.710 4.310 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.730 0.840 9.100 1.210 ;
        RECT  8.730 0.330 9.010 2.100 ;
        RECT  8.660 0.330 9.010 0.830 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.690 3.530 9.100 3.960 ;
        RECT  8.690 2.740 8.970 4.470 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.000 1.280 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.170 1.500 8.450 3.330 ;
        RECT  7.210 2.260 7.410 3.000 ;
        RECT  5.320 1.680 5.600 2.540 ;
        RECT  3.030 1.770 3.310 2.540 ;
        RECT  2.970 2.260 3.270 3.050 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.050 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.170 -0.140 8.450 0.610 ;
        RECT  5.080 -0.140 5.350 0.560 ;
        RECT  2.500 -0.140 2.780 0.320 ;
        RECT  0.000 4.660 9.200 4.940 ;
        RECT  8.210 4.020 8.450 4.940 ;
        RECT  7.130 4.300 7.410 4.940 ;
        RECT  4.770 4.480 5.050 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.210 1.030 3.380 ;
        RECT  0.870 3.210 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.050 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.640 1.130 2.560 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.640 1.130 1.800 1.820 ;
        RECT  0.100 1.660 1.800 1.820 ;
        RECT  1.070 0.300 2.240 0.460 ;
        RECT  2.070 0.300 2.240 0.640 ;
        RECT  3.100 0.320 3.380 0.640 ;
        RECT  2.070 0.480 3.380 0.640 ;
        RECT  1.070 0.300 1.310 0.830 ;
        RECT  1.570 0.620 1.850 0.960 ;
        RECT  3.580 0.340 3.860 0.960 ;
        RECT  1.570 0.800 3.860 0.960 ;
        RECT  3.610 2.700 3.970 2.960 ;
        RECT  3.610 2.700 3.790 4.160 ;
        RECT  3.350 3.940 3.790 4.160 ;
        RECT  2.710 1.410 4.010 1.610 ;
        RECT  2.070 1.600 2.870 1.770 ;
        RECT  4.090 0.340 4.560 0.670 ;
        RECT  4.240 0.340 4.560 1.200 ;
        RECT  4.240 1.040 5.770 1.200 ;
        RECT  4.240 0.340 4.480 1.650 ;
        RECT  4.770 3.020 5.920 3.180 ;
        RECT  5.610 3.020 5.920 3.720 ;
        RECT  4.770 3.020 4.930 3.660 ;
        RECT  4.590 3.440 4.930 3.660 ;
        RECT  5.610 3.430 6.000 3.720 ;
        RECT  5.610 3.020 5.850 4.150 ;
        RECT  5.560 3.900 5.850 4.150 ;
        RECT  4.190 2.700 6.670 2.860 ;
        RECT  4.190 2.700 4.350 3.360 ;
        RECT  3.950 3.120 4.230 4.150 ;
        RECT  5.930 1.040 6.900 1.320 ;
        RECT  5.930 1.040 6.090 1.520 ;
        RECT  4.810 1.360 6.090 1.520 ;
        RECT  4.810 1.360 4.970 2.040 ;
        RECT  3.480 1.810 4.970 2.040 ;
        RECT  5.600 0.460 5.880 0.880 ;
        RECT  6.200 0.340 6.480 0.880 ;
        RECT  4.720 0.720 7.230 0.880 ;
        RECT  7.070 0.720 7.230 1.640 ;
        RECT  6.700 1.480 7.230 1.640 ;
        RECT  5.800 1.680 6.880 1.840 ;
        RECT  6.700 1.480 6.880 1.860 ;
        RECT  6.530 1.660 6.880 1.860 ;
        RECT  6.130 3.080 6.410 3.300 ;
        RECT  6.160 3.160 7.430 3.320 ;
        RECT  7.270 3.160 7.430 3.750 ;
        RECT  7.270 3.500 7.610 3.750 ;
        RECT  6.160 3.160 6.440 4.180 ;
        RECT  6.100 3.900 6.440 4.180 ;
        RECT  7.730 2.700 7.930 3.390 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  7.770 3.510 8.450 3.790 ;
        RECT  6.760 3.510 7.110 4.070 ;
        RECT  6.760 3.910 7.930 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.450 4.160 5.370 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.210 4.160 5.370 4.500 ;
        RECT  7.770 2.700 7.930 4.490 ;
        RECT  7.650 3.910 7.930 4.490 ;
        RECT  4.450 4.160 4.610 4.500 ;
        RECT  3.030 4.340 4.610 4.500 ;
        RECT  6.760 3.510 6.920 4.500 ;
        RECT  5.210 4.340 6.920 4.500 ;
        RECT  6.800 0.340 7.550 0.500 ;
        RECT  7.390 1.030 8.510 1.250 ;
        RECT  7.390 0.340 7.550 1.960 ;
        RECT  7.040 1.800 7.550 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.200 3.540 ;
        RECT  3.460 1.070 7.540 3.600 ;
        RECT  2.860 1.140 9.200 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.330 1.140 9.200 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.330 4.800 ;
        RECT  0.000 3.660 9.200 4.800 ;
        RECT  0.000 0.000 9.200 1.070 ;
        RECT  0.000 0.000 3.460 1.140 ;
        RECT  7.540 0.000 9.200 1.140 ;
    END
END SDFEM2HM

MACRO SDFEM1HM
    CLASS CORE ;
    FOREIGN SDFEM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.635  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.250 3.420 5.450 3.620 ;
        LAYER ME2 ;
        RECT  5.250 3.240 5.500 3.960 ;
        LAYER ME1 ;
        RECT  5.130 3.340 5.450 3.750 ;
        RECT  5.130 3.340 5.400 4.000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.230 3.220 1.610 3.680 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.150  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.540 0.710 4.310 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.800 0.840 9.100 1.210 ;
        RECT  8.800 0.330 9.010 1.760 ;
        RECT  8.730 0.330 9.010 0.830 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.760 3.530 9.100 3.960 ;
        RECT  8.760 2.940 9.040 4.470 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 3.240 3.430 3.780 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.630 1.000 1.280 1.500 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.240 1.500 8.520 3.330 ;
        RECT  7.210 2.260 7.410 3.000 ;
        RECT  5.360 1.680 5.640 2.540 ;
        RECT  3.070 1.770 3.350 2.540 ;
        RECT  2.970 2.260 3.270 3.050 ;
        RECT  0.660 1.980 0.940 2.540 ;
        RECT  0.620 2.260 0.910 3.050 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.240 -0.140 8.520 0.610 ;
        RECT  5.120 -0.140 5.390 0.560 ;
        RECT  2.540 -0.140 2.820 0.320 ;
        RECT  0.000 4.660 9.200 4.940 ;
        RECT  8.280 4.190 8.520 4.940 ;
        RECT  7.130 4.300 7.410 4.940 ;
        RECT  4.770 4.480 5.050 4.940 ;
        RECT  2.590 4.470 2.870 4.940 ;
        RECT  0.660 4.470 0.940 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 3.210 1.030 3.380 ;
        RECT  0.870 3.210 1.030 4.180 ;
        RECT  0.870 4.020 1.370 4.180 ;
        RECT  1.210 4.020 1.370 4.500 ;
        RECT  0.140 2.880 0.340 4.470 ;
        RECT  1.210 4.340 2.190 4.500 ;
        RECT  1.430 2.700 2.510 2.910 ;
        RECT  1.430 2.700 1.990 3.050 ;
        RECT  1.800 2.700 1.990 4.180 ;
        RECT  1.610 3.920 1.990 4.180 ;
        RECT  1.680 1.130 2.600 1.350 ;
        RECT  0.100 0.310 0.380 1.820 ;
        RECT  1.680 1.130 1.840 1.820 ;
        RECT  0.100 1.660 1.840 1.820 ;
        RECT  1.070 0.300 2.280 0.460 ;
        RECT  2.110 0.300 2.280 0.640 ;
        RECT  3.140 0.320 3.420 0.640 ;
        RECT  2.110 0.480 3.420 0.640 ;
        RECT  1.070 0.300 1.310 0.830 ;
        RECT  1.610 0.620 1.890 0.960 ;
        RECT  3.620 0.340 3.900 0.960 ;
        RECT  1.610 0.800 3.900 0.960 ;
        RECT  3.670 2.700 3.970 2.960 ;
        RECT  3.670 2.700 3.850 4.160 ;
        RECT  3.350 3.940 3.850 4.160 ;
        RECT  2.750 1.410 4.050 1.610 ;
        RECT  2.110 1.600 2.910 1.770 ;
        RECT  4.130 0.340 4.460 0.670 ;
        RECT  4.280 0.340 4.460 1.650 ;
        RECT  4.280 1.040 5.810 1.200 ;
        RECT  4.280 1.040 4.560 1.650 ;
        RECT  4.770 3.020 5.920 3.180 ;
        RECT  5.610 3.020 5.920 3.720 ;
        RECT  4.770 3.020 4.930 3.660 ;
        RECT  4.590 3.440 4.930 3.660 ;
        RECT  5.610 3.430 6.000 3.720 ;
        RECT  5.610 3.020 5.850 4.150 ;
        RECT  5.560 3.900 5.850 4.150 ;
        RECT  4.190 2.700 6.670 2.860 ;
        RECT  4.190 2.700 4.350 3.400 ;
        RECT  4.010 3.120 4.290 4.150 ;
        RECT  5.970 1.040 6.940 1.320 ;
        RECT  5.970 1.040 6.130 1.520 ;
        RECT  4.850 1.360 6.130 1.520 ;
        RECT  4.850 1.360 5.010 2.040 ;
        RECT  3.520 1.810 5.010 2.040 ;
        RECT  5.640 0.460 5.920 0.880 ;
        RECT  6.240 0.340 6.520 0.880 ;
        RECT  4.760 0.720 7.270 0.880 ;
        RECT  7.110 0.720 7.270 1.640 ;
        RECT  6.740 1.480 7.270 1.640 ;
        RECT  5.840 1.680 6.920 1.840 ;
        RECT  6.740 1.480 6.920 1.860 ;
        RECT  6.570 1.660 6.920 1.860 ;
        RECT  6.130 3.080 6.410 3.300 ;
        RECT  6.160 3.160 7.430 3.320 ;
        RECT  7.270 3.160 7.430 3.750 ;
        RECT  7.270 3.500 7.610 3.750 ;
        RECT  6.160 3.160 6.440 4.180 ;
        RECT  6.100 3.900 6.440 4.180 ;
        RECT  7.730 2.700 7.930 3.390 ;
        RECT  7.770 2.700 7.930 4.490 ;
        RECT  2.330 3.360 2.660 3.640 ;
        RECT  7.770 3.510 8.520 3.790 ;
        RECT  6.760 3.510 7.110 4.070 ;
        RECT  6.760 3.910 8.010 4.070 ;
        RECT  2.500 3.360 2.660 4.250 ;
        RECT  2.500 4.090 3.190 4.250 ;
        RECT  4.450 4.160 5.370 4.320 ;
        RECT  3.030 4.090 3.190 4.500 ;
        RECT  5.210 4.160 5.370 4.500 ;
        RECT  7.770 3.510 8.010 4.490 ;
        RECT  7.730 3.910 8.010 4.490 ;
        RECT  4.450 4.160 4.610 4.500 ;
        RECT  3.030 4.340 4.610 4.500 ;
        RECT  6.760 3.510 6.920 4.500 ;
        RECT  5.210 4.340 6.920 4.500 ;
        RECT  6.840 0.340 7.590 0.500 ;
        RECT  7.430 1.030 8.580 1.250 ;
        RECT  7.430 0.340 7.590 1.960 ;
        RECT  7.080 1.800 7.590 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.200 3.540 ;
        RECT  3.500 1.070 7.580 3.600 ;
        RECT  2.860 1.140 9.200 3.600 ;
        RECT  0.000 1.140 1.170 3.660 ;
        RECT  6.330 1.140 9.200 3.660 ;
        LAYER VTNH ;
        RECT  1.170 3.540 2.860 4.800 ;
        RECT  1.170 3.600 6.330 4.800 ;
        RECT  0.000 3.660 9.200 4.800 ;
        RECT  0.000 0.000 9.200 1.070 ;
        RECT  0.000 0.000 3.500 1.140 ;
        RECT  7.580 0.000 9.200 1.140 ;
    END
END SDFEM1HM

MACRO SDFCRSM8HM
    CLASS CORE ;
    FOREIGN SDFCRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.383  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.580 1.280 2.780 1.480 ;
        LAYER ME2 ;
        RECT  2.500 1.170 2.780 1.560 ;
        LAYER ME1 ;
        RECT  2.580 1.040 2.950 1.560 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER ME1  ;
        ANTENNAGATEAREA 0.245  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.806  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  15.300 1.020 15.500 1.220 ;
        LAYER ME2 ;
        RECT  15.300 0.810 15.500 1.560 ;
        LAYER ME1 ;
        RECT  15.030 0.940 15.600 1.220 ;
        END
    END RB
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.270 1.300 18.750 1.600 ;
        RECT  18.370 0.300 18.610 1.600 ;
        RECT  17.270 0.300 17.500 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  20.680 0.300 20.960 2.080 ;
        RECT  19.640 0.840 20.960 1.160 ;
        RECT  19.640 0.300 19.920 1.160 ;
        RECT  19.640 0.300 19.910 2.080 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.052  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 21.600 2.540 ;
        RECT  21.200 1.500 21.480 2.540 ;
        RECT  20.160 1.500 20.440 2.540 ;
        RECT  19.080 2.080 19.360 2.540 ;
        RECT  17.870 2.080 18.150 2.540 ;
        RECT  16.590 2.080 16.870 2.540 ;
        RECT  15.390 2.080 15.670 2.540 ;
        RECT  13.830 1.820 14.030 2.540 ;
        RECT  12.230 2.080 12.510 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 21.600 0.140 ;
        RECT  21.200 -0.140 21.480 0.580 ;
        RECT  20.160 -0.140 20.440 0.580 ;
        RECT  19.120 -0.140 19.400 0.580 ;
        RECT  17.760 -0.140 18.040 0.590 ;
        RECT  16.580 -0.140 16.860 0.320 ;
        RECT  13.920 -0.140 14.200 0.540 ;
        RECT  12.050 -0.140 12.330 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.620 0.880 ;
        RECT  1.460 0.880 1.660 1.230 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.540 0.840 ;
        RECT  2.180 0.620 2.380 1.780 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.680 1.480 1.880 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.680 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.780 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  1.780 0.300 1.980 0.680 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.050 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.050 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  16.090 1.240 16.410 1.600 ;
        RECT  13.510 1.390 16.410 1.600 ;
        RECT  11.910 1.760 12.910 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.730 1.760 12.910 2.100 ;
        RECT  11.910 1.760 12.070 2.100 ;
        RECT  10.540 1.940 12.070 2.100 ;
        RECT  13.510 1.390 13.670 2.100 ;
        RECT  12.730 1.940 13.670 2.100 ;
        RECT  14.680 0.620 15.930 0.780 ;
        RECT  15.770 0.620 15.930 0.960 ;
        RECT  15.770 0.800 16.790 0.960 ;
        RECT  14.680 0.620 14.840 1.180 ;
        RECT  11.910 1.020 14.840 1.180 ;
        RECT  16.630 0.800 16.790 1.920 ;
        RECT  14.310 1.760 16.790 1.920 ;
        RECT  14.310 1.760 14.660 2.100 ;
        RECT  14.360 0.300 16.250 0.460 ;
        RECT  16.090 0.300 16.250 0.640 ;
        RECT  16.090 0.480 17.110 0.640 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.990 0.540 13.270 0.860 ;
        RECT  14.360 0.300 14.520 0.860 ;
        RECT  11.460 0.700 14.520 0.860 ;
        RECT  19.180 1.060 19.460 1.340 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.350 1.600 ;
        RECT  16.950 0.480 17.110 1.920 ;
        RECT  13.070 1.440 13.350 1.780 ;
        RECT  19.180 1.060 19.340 1.920 ;
        RECT  16.950 1.760 19.340 1.920 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.980 2.400 ;
        RECT  17.080 1.080 18.930 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 21.600 2.400 ;
        RECT  11.090 1.140 21.600 2.400 ;
        RECT  0.000 1.210 21.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 21.600 1.070 ;
        RECT  11.980 0.000 21.600 1.080 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.980 0.000 17.080 1.140 ;
        RECT  18.930 0.000 21.600 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCRSM8HM

MACRO SDFCRSM4HM
    CLASS CORE ;
    FOREIGN SDFCRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.973  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  15.030 1.280 15.230 1.480 ;
        LAYER ME2 ;
        RECT  14.900 1.220 15.230 1.560 ;
        LAYER ME1 ;
        RECT  15.030 0.940 15.350 1.560 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.110  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.580 1.280 2.780 1.480 ;
        LAYER ME2 ;
        RECT  2.500 1.170 2.780 1.560 ;
        LAYER ME1 ;
        RECT  2.580 1.040 2.950 1.560 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.611  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.500 1.200 16.930 1.600 ;
        RECT  16.610 0.300 16.930 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.770 0.840 18.300 1.160 ;
        RECT  17.770 0.840 18.110 2.080 ;
        RECT  17.770 0.300 18.070 2.080 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.800 2.540 ;
        RECT  18.310 1.500 18.590 2.540 ;
        RECT  17.230 2.080 17.510 2.540 ;
        RECT  15.390 2.080 15.670 2.540 ;
        RECT  13.830 1.820 14.030 2.540 ;
        RECT  12.230 2.080 12.510 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.800 0.140 ;
        RECT  18.310 -0.140 18.590 0.580 ;
        RECT  17.270 -0.140 17.550 0.580 ;
        RECT  16.150 -0.140 16.430 0.590 ;
        RECT  13.920 -0.140 14.200 0.540 ;
        RECT  12.050 -0.140 12.330 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.620 0.880 ;
        RECT  1.460 0.880 1.660 1.230 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.540 0.840 ;
        RECT  2.180 0.620 2.380 1.780 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.680 1.480 1.880 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.680 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.780 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  1.780 0.300 1.980 0.680 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.050 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.050 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  13.510 1.390 14.870 1.600 ;
        RECT  11.910 1.760 12.910 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.730 1.760 12.910 2.100 ;
        RECT  11.910 1.760 12.070 2.100 ;
        RECT  10.540 1.940 12.070 2.100 ;
        RECT  13.510 1.390 13.670 2.100 ;
        RECT  12.730 1.940 13.670 2.100 ;
        RECT  14.680 0.620 15.670 0.780 ;
        RECT  14.680 0.620 14.840 1.180 ;
        RECT  11.910 1.020 14.840 1.180 ;
        RECT  15.510 0.620 15.670 1.920 ;
        RECT  14.310 1.760 15.670 1.920 ;
        RECT  14.310 1.760 14.660 2.100 ;
        RECT  14.360 0.300 15.990 0.460 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.990 0.540 13.270 0.860 ;
        RECT  14.360 0.300 14.520 0.860 ;
        RECT  11.460 0.700 14.520 0.860 ;
        RECT  17.330 1.060 17.610 1.340 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.350 1.600 ;
        RECT  15.830 0.300 15.990 1.920 ;
        RECT  13.070 1.440 13.350 1.780 ;
        RECT  17.330 1.060 17.490 1.920 ;
        RECT  15.830 1.760 17.490 1.920 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.980 2.400 ;
        RECT  15.830 1.080 17.120 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 18.800 2.400 ;
        RECT  11.090 1.140 18.800 2.400 ;
        RECT  0.000 1.210 18.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.800 1.070 ;
        RECT  11.980 0.000 18.800 1.080 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.980 0.000 15.830 1.140 ;
        RECT  17.120 0.000 18.800 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCRSM4HM

MACRO SDFCRSM2HM
    CLASS CORE ;
    FOREIGN SDFCRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.110  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.580 1.280 2.780 1.480 ;
        LAYER ME2 ;
        RECT  2.500 1.120 2.780 1.560 ;
        LAYER ME1 ;
        RECT  2.580 1.040 2.950 1.560 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.783  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  14.980 1.280 15.180 1.480 ;
        LAYER ME2 ;
        RECT  14.900 1.170 15.180 1.560 ;
        LAYER ME1 ;
        RECT  14.980 0.940 15.240 1.560 ;
        END
    END RB
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.040 0.300 16.340 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.180 0.300 17.500 2.080 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.600 2.540 ;
        RECT  16.640 2.080 16.920 2.540 ;
        RECT  15.340 2.080 15.620 2.540 ;
        RECT  13.780 1.820 13.980 2.540 ;
        RECT  12.180 2.080 12.460 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.600 0.140 ;
        RECT  16.680 -0.140 16.960 0.580 ;
        RECT  13.870 -0.140 14.150 0.540 ;
        RECT  12.000 -0.140 12.280 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.620 0.880 ;
        RECT  1.460 0.870 1.660 1.230 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.540 0.840 ;
        RECT  2.180 0.620 2.380 1.780 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.680 1.480 1.880 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.680 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.780 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  1.780 0.300 1.980 0.680 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.060 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.060 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  13.460 1.390 14.820 1.600 ;
        RECT  11.860 1.760 12.860 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.680 1.760 12.860 2.100 ;
        RECT  11.860 1.760 12.020 2.100 ;
        RECT  10.540 1.940 12.020 2.100 ;
        RECT  13.460 1.390 13.620 2.100 ;
        RECT  12.680 1.940 13.620 2.100 ;
        RECT  14.630 0.620 15.560 0.780 ;
        RECT  14.630 0.620 14.790 1.220 ;
        RECT  11.900 1.020 14.790 1.220 ;
        RECT  15.400 0.620 15.560 1.920 ;
        RECT  14.260 1.760 15.560 1.920 ;
        RECT  14.260 1.760 14.610 2.100 ;
        RECT  14.310 0.300 15.880 0.460 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.940 0.540 13.220 0.860 ;
        RECT  14.310 0.300 14.470 0.860 ;
        RECT  11.460 0.700 14.470 0.860 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.300 1.600 ;
        RECT  15.720 0.300 15.880 1.920 ;
        RECT  13.020 1.440 13.300 1.780 ;
        RECT  16.740 1.060 17.020 1.920 ;
        RECT  15.720 1.760 17.020 1.920 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.940 2.400 ;
        RECT  15.720 1.080 16.610 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 17.600 2.400 ;
        RECT  11.090 1.140 17.600 2.400 ;
        RECT  0.000 1.210 17.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.600 1.070 ;
        RECT  11.940 0.000 17.600 1.080 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.940 0.000 15.720 1.140 ;
        RECT  16.610 0.000 17.600 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCRSM2HM

MACRO SDFCRSM1HM
    CLASS CORE ;
    FOREIGN SDFCRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        ANTENNAGATEAREA 0.102  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.569  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.880 1.100 2.080 1.300 ;
        LAYER ME2 ;
        RECT  1.700 0.840 2.080 1.380 ;
        LAYER ME1 ;
        RECT  1.820 1.040 2.180 1.380 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.783  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  14.980 1.280 15.180 1.480 ;
        LAYER ME2 ;
        RECT  14.900 1.170 15.180 1.560 ;
        LAYER ME1 ;
        RECT  14.980 0.940 15.240 1.560 ;
        END
    END RB
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.332  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.040 0.300 16.340 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.180 0.300 17.500 1.800 ;
        END
    END QB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.600 2.540 ;
        RECT  16.640 2.080 16.920 2.540 ;
        RECT  15.340 2.080 15.620 2.540 ;
        RECT  13.780 1.820 13.980 2.540 ;
        RECT  12.180 2.080 12.460 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.600 0.140 ;
        RECT  16.680 -0.140 16.960 0.580 ;
        RECT  13.870 -0.140 14.150 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 2.540 0.880 ;
        RECT  2.350 0.720 2.540 1.220 ;
        RECT  2.350 0.940 2.770 1.220 ;
        RECT  1.460 0.720 1.660 1.270 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.640 1.540 1.920 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.640 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.740 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  1.740 0.300 2.060 0.540 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.060 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.060 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  13.460 1.390 14.820 1.600 ;
        RECT  11.860 1.760 12.860 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.680 1.760 12.860 2.100 ;
        RECT  11.860 1.760 12.020 2.100 ;
        RECT  10.540 1.940 12.020 2.100 ;
        RECT  13.460 1.390 13.620 2.100 ;
        RECT  12.680 1.940 13.620 2.100 ;
        RECT  14.630 0.620 15.560 0.780 ;
        RECT  14.630 0.620 14.790 1.220 ;
        RECT  11.900 1.020 14.790 1.220 ;
        RECT  15.400 0.620 15.560 1.920 ;
        RECT  14.260 1.760 15.560 1.920 ;
        RECT  14.260 1.760 14.610 2.100 ;
        RECT  14.310 0.300 15.880 0.460 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.420 0.540 12.700 0.860 ;
        RECT  14.310 0.300 14.470 0.860 ;
        RECT  11.460 0.700 14.470 0.860 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.300 1.600 ;
        RECT  15.720 0.300 15.880 1.920 ;
        RECT  13.020 1.440 13.300 1.780 ;
        RECT  16.740 1.060 17.020 1.920 ;
        RECT  15.720 1.760 17.020 1.920 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.940 2.400 ;
        RECT  15.720 1.080 16.610 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 17.600 2.400 ;
        RECT  11.090 1.140 17.600 2.400 ;
        RECT  0.000 1.210 17.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.600 1.070 ;
        RECT  11.940 0.000 17.600 1.080 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.940 0.000 15.720 1.140 ;
        RECT  16.610 0.000 17.600 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCRSM1HM

MACRO SDFCQRSM8HM
    CLASS CORE ;
    FOREIGN SDFCQRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.383  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.580 1.280 2.780 1.480 ;
        LAYER ME2 ;
        RECT  2.500 1.170 2.780 1.560 ;
        LAYER ME1 ;
        RECT  2.580 1.040 2.950 1.560 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER ME1  ;
        ANTENNAGATEAREA 0.245  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.806  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  15.300 1.020 15.500 1.220 ;
        LAYER ME2 ;
        RECT  15.300 0.810 15.500 1.560 ;
        LAYER ME1 ;
        RECT  15.030 0.940 15.600 1.220 ;
        END
    END RB
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  18.180 1.300 18.490 2.070 ;
        RECT  18.210 0.300 18.490 2.070 ;
        RECT  17.150 1.300 18.490 1.660 ;
        RECT  17.150 1.300 17.440 2.100 ;
        RECT  17.150 0.300 17.410 2.100 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.052  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 19.200 2.540 ;
        RECT  18.710 1.390 18.990 2.540 ;
        RECT  17.670 1.890 17.950 2.540 ;
        RECT  16.590 2.080 16.870 2.540 ;
        RECT  15.390 2.080 15.670 2.540 ;
        RECT  13.830 1.820 14.030 2.540 ;
        RECT  12.230 2.080 12.510 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 19.200 0.140 ;
        RECT  18.710 -0.140 18.990 0.580 ;
        RECT  17.670 -0.140 17.950 0.670 ;
        RECT  16.080 -0.140 16.920 0.550 ;
        RECT  13.920 -0.140 14.200 0.540 ;
        RECT  12.050 -0.140 12.330 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.620 0.880 ;
        RECT  1.460 0.880 1.660 1.230 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.540 0.840 ;
        RECT  2.180 0.620 2.380 1.780 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.680 1.480 1.880 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.680 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.780 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  1.780 0.300 1.980 0.680 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.050 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.050 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.990 0.540 13.270 0.860 ;
        RECT  11.460 0.700 13.350 0.860 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.350 1.600 ;
        RECT  13.070 1.440 13.350 1.780 ;
        RECT  16.090 1.240 16.410 1.600 ;
        RECT  13.510 1.390 16.410 1.600 ;
        RECT  11.910 1.760 12.910 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.730 1.760 12.910 2.100 ;
        RECT  11.910 1.760 12.070 2.100 ;
        RECT  10.540 1.940 12.070 2.100 ;
        RECT  13.510 1.390 13.670 2.100 ;
        RECT  12.730 1.940 13.670 2.100 ;
        RECT  14.680 0.620 15.930 0.780 ;
        RECT  15.770 0.620 15.930 0.960 ;
        RECT  15.770 0.800 16.790 0.960 ;
        RECT  14.680 0.620 14.840 1.180 ;
        RECT  11.910 1.020 14.840 1.180 ;
        RECT  16.630 0.800 16.790 1.920 ;
        RECT  14.310 1.760 16.790 1.920 ;
        RECT  14.310 1.760 14.660 2.100 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.980 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 19.200 2.400 ;
        RECT  11.090 1.140 19.200 2.400 ;
        RECT  0.000 1.210 19.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 19.200 1.070 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.980 0.000 19.200 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCQRSM8HM

MACRO SDFCQRSM4HM
    CLASS CORE ;
    FOREIGN SDFCQRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.783  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  15.030 1.280 15.230 1.480 ;
        LAYER ME2 ;
        RECT  14.900 1.220 15.230 1.560 ;
        LAYER ME1 ;
        RECT  15.030 0.940 15.290 1.560 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.110  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.580 1.280 2.780 1.480 ;
        LAYER ME2 ;
        RECT  2.500 1.170 2.780 1.560 ;
        LAYER ME1 ;
        RECT  2.580 1.040 2.950 1.560 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.100 1.200 16.510 2.100 ;
        RECT  16.170 0.300 16.510 2.100 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.200 2.540 ;
        RECT  16.750 1.400 17.030 2.540 ;
        RECT  15.770 1.410 15.930 2.540 ;
        RECT  13.830 1.820 14.030 2.540 ;
        RECT  12.230 2.080 12.510 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.200 0.140 ;
        RECT  16.750 -0.140 17.030 0.580 ;
        RECT  15.770 -0.140 15.990 0.710 ;
        RECT  13.920 -0.140 14.200 0.540 ;
        RECT  12.050 -0.140 12.330 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.620 0.880 ;
        RECT  1.460 0.880 1.660 1.230 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.540 0.840 ;
        RECT  2.180 0.620 2.380 1.780 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.680 1.480 1.880 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.680 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.780 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  1.780 0.300 1.980 0.680 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.050 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.050 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.990 0.540 13.270 0.860 ;
        RECT  11.460 0.700 13.270 0.860 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.350 1.600 ;
        RECT  13.070 1.440 13.350 1.780 ;
        RECT  13.510 1.390 14.870 1.600 ;
        RECT  11.910 1.760 12.910 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.730 1.760 12.910 2.100 ;
        RECT  11.910 1.760 12.070 2.100 ;
        RECT  10.540 1.940 12.070 2.100 ;
        RECT  13.510 1.390 13.670 2.100 ;
        RECT  12.730 1.940 13.670 2.100 ;
        RECT  14.680 0.620 15.610 0.780 ;
        RECT  14.680 0.620 14.840 1.180 ;
        RECT  11.910 1.020 14.840 1.180 ;
        RECT  15.450 0.970 15.830 1.250 ;
        RECT  15.450 0.620 15.610 1.920 ;
        RECT  14.310 1.760 15.610 1.920 ;
        RECT  14.310 1.760 14.660 2.100 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.980 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 17.200 2.400 ;
        RECT  11.090 1.140 17.200 2.400 ;
        RECT  0.000 1.210 17.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.200 1.070 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.980 0.000 17.200 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCQRSM4HM

MACRO SDFCQRSM2HM
    CLASS CORE ;
    FOREIGN SDFCQRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.110  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.580 1.280 2.780 1.480 ;
        LAYER ME2 ;
        RECT  2.500 1.120 2.780 1.560 ;
        LAYER ME1 ;
        RECT  2.580 1.040 2.950 1.560 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.783  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  14.980 1.280 15.180 1.480 ;
        LAYER ME2 ;
        RECT  14.900 1.170 15.180 1.560 ;
        LAYER ME1 ;
        RECT  14.980 0.940 15.240 1.560 ;
        END
    END RB
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.780 0.840 16.360 1.160 ;
        RECT  15.780 0.300 16.140 2.100 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.800 2.540 ;
        RECT  16.340 1.440 16.620 2.540 ;
        RECT  15.340 2.080 15.620 2.540 ;
        RECT  13.780 1.820 13.980 2.540 ;
        RECT  12.180 2.080 12.460 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.800 0.140 ;
        RECT  16.340 -0.140 16.620 0.580 ;
        RECT  13.870 -0.140 14.150 0.540 ;
        RECT  12.000 -0.140 12.280 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.620 0.880 ;
        RECT  1.460 0.870 1.660 1.230 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.540 0.840 ;
        RECT  2.180 0.620 2.380 1.780 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.680 1.480 1.880 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.680 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.780 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  1.780 0.300 1.980 0.680 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.060 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.060 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.940 0.540 13.220 0.860 ;
        RECT  11.460 0.700 13.220 0.860 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.300 1.600 ;
        RECT  13.020 1.440 13.300 1.780 ;
        RECT  13.460 1.390 14.820 1.600 ;
        RECT  11.860 1.760 12.860 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.680 1.760 12.860 2.100 ;
        RECT  11.860 1.760 12.020 2.100 ;
        RECT  10.540 1.940 12.020 2.100 ;
        RECT  13.460 1.390 13.620 2.100 ;
        RECT  12.680 1.940 13.620 2.100 ;
        RECT  14.630 0.620 15.560 0.780 ;
        RECT  14.630 0.620 14.790 1.220 ;
        RECT  11.900 1.020 14.790 1.220 ;
        RECT  15.400 0.620 15.560 1.920 ;
        RECT  14.260 1.760 15.560 1.920 ;
        RECT  14.260 1.760 14.610 2.100 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.940 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 16.800 2.400 ;
        RECT  11.090 1.140 16.800 2.400 ;
        RECT  0.000 1.210 16.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.800 1.070 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.940 0.000 16.800 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCQRSM2HM

MACRO SDFCQRSM1HM
    CLASS CORE ;
    FOREIGN SDFCQRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        ANTENNAGATEAREA 0.102  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.569  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.880 1.100 2.080 1.300 ;
        LAYER ME2 ;
        RECT  1.700 0.840 2.080 1.380 ;
        LAYER ME1 ;
        RECT  1.820 1.040 2.180 1.380 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.783  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  14.980 1.280 15.180 1.480 ;
        LAYER ME2 ;
        RECT  14.900 1.170 15.180 1.560 ;
        LAYER ME1 ;
        RECT  14.980 0.940 15.240 1.560 ;
        END
    END RB
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.150 1.040 3.500 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.820 0.840 16.300 1.160 ;
        RECT  15.820 0.300 16.120 1.770 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 1.830 10.320 2.100 ;
        RECT  9.700 1.170 9.900 2.100 ;
        RECT  9.200 1.170 9.900 1.340 ;
        RECT  9.200 0.980 9.450 1.340 ;
        END
    END SB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.800 2.540 ;
        RECT  16.340 1.570 16.620 2.540 ;
        RECT  15.340 2.080 15.620 2.540 ;
        RECT  13.780 1.820 13.980 2.540 ;
        RECT  12.180 2.080 12.460 2.540 ;
        RECT  8.560 1.860 8.840 2.540 ;
        RECT  6.840 1.440 7.120 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.800 0.140 ;
        RECT  16.340 -0.140 16.620 0.580 ;
        RECT  13.870 -0.140 14.150 0.540 ;
        RECT  8.240 -0.140 8.400 0.640 ;
        RECT  4.420 -0.140 4.580 0.420 ;
        RECT  3.020 -0.140 3.180 0.420 ;
        RECT  0.660 -0.140 0.940 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 2.540 0.880 ;
        RECT  2.350 0.720 2.540 1.220 ;
        RECT  2.350 0.940 2.770 1.220 ;
        RECT  1.460 0.720 1.660 1.270 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  3.660 0.900 4.760 1.180 ;
        RECT  3.660 0.620 3.940 1.660 ;
        RECT  5.060 0.620 5.340 1.660 ;
        RECT  4.540 1.500 5.340 1.660 ;
        RECT  2.540 1.760 3.500 1.920 ;
        RECT  1.640 1.540 1.920 2.100 ;
        RECT  3.340 1.760 3.500 2.100 ;
        RECT  2.540 1.760 2.700 2.100 ;
        RECT  1.640 1.940 2.700 2.100 ;
        RECT  5.060 1.860 5.380 2.100 ;
        RECT  3.340 1.940 5.380 2.100 ;
        RECT  1.740 0.300 2.860 0.460 ;
        RECT  3.340 0.300 4.260 0.460 ;
        RECT  4.740 0.300 5.820 0.460 ;
        RECT  1.740 0.300 2.060 0.540 ;
        RECT  2.700 0.300 2.860 0.740 ;
        RECT  4.100 0.300 4.260 0.740 ;
        RECT  3.340 0.300 3.500 0.740 ;
        RECT  2.700 0.580 3.500 0.740 ;
        RECT  4.740 0.300 4.900 0.740 ;
        RECT  4.100 0.580 4.900 0.740 ;
        RECT  5.540 0.300 5.820 0.880 ;
        RECT  6.060 0.620 7.760 0.780 ;
        RECT  7.600 0.620 7.760 1.280 ;
        RECT  7.600 1.120 8.680 1.280 ;
        RECT  6.060 0.620 6.220 1.360 ;
        RECT  5.580 1.200 6.220 1.360 ;
        RECT  5.580 1.200 5.860 2.080 ;
        RECT  8.880 0.620 9.450 0.820 ;
        RECT  6.830 1.080 7.440 1.280 ;
        RECT  7.280 1.080 7.440 1.700 ;
        RECT  8.880 0.620 9.040 1.700 ;
        RECT  7.280 1.540 9.400 1.700 ;
        RECT  9.080 1.540 9.400 1.740 ;
        RECT  7.920 1.540 8.200 1.760 ;
        RECT  6.480 0.300 8.080 0.460 ;
        RECT  8.560 0.300 11.300 0.460 ;
        RECT  7.920 0.300 8.080 0.960 ;
        RECT  8.560 0.300 8.720 0.960 ;
        RECT  7.920 0.800 8.720 0.960 ;
        RECT  9.620 0.300 9.900 0.990 ;
        RECT  11.140 0.300 11.300 1.660 ;
        RECT  11.460 0.490 11.790 0.860 ;
        RECT  12.420 0.540 12.700 0.860 ;
        RECT  11.460 0.700 12.700 0.860 ;
        RECT  11.460 0.490 11.740 1.600 ;
        RECT  11.460 1.440 13.300 1.600 ;
        RECT  13.020 1.440 13.300 1.780 ;
        RECT  13.460 1.390 14.820 1.600 ;
        RECT  11.860 1.760 12.860 1.920 ;
        RECT  10.540 0.620 10.820 2.100 ;
        RECT  12.680 1.760 12.860 2.100 ;
        RECT  11.860 1.760 12.020 2.100 ;
        RECT  10.540 1.940 12.020 2.100 ;
        RECT  13.460 1.390 13.620 2.100 ;
        RECT  12.680 1.940 13.620 2.100 ;
        RECT  14.630 0.620 15.560 0.780 ;
        RECT  14.630 0.620 14.790 1.220 ;
        RECT  11.900 1.020 14.790 1.220 ;
        RECT  15.400 0.620 15.560 1.920 ;
        RECT  14.260 1.760 15.560 1.920 ;
        RECT  14.260 1.760 14.610 2.100 ;
        LAYER VTPH ;
        RECT  11.090 1.070 11.940 2.400 ;
        RECT  0.000 1.140 7.920 2.400 ;
        RECT  9.600 1.170 16.800 2.400 ;
        RECT  11.090 1.140 16.800 2.400 ;
        RECT  0.000 1.210 16.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.800 1.070 ;
        RECT  0.000 0.000 11.090 1.140 ;
        RECT  11.940 0.000 16.800 1.140 ;
        RECT  7.920 0.000 11.090 1.170 ;
        RECT  7.920 0.000 9.600 1.210 ;
    END
END SDFCQRSM1HM

MACRO SDFCQM8HM
    CLASS CORE ;
    FOREIGN SDFCQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.060 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.060 3.100 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.039  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.810 0.840 14.090 2.100 ;
        RECT  13.870 0.460 14.090 2.100 ;
        RECT  12.750 0.840 14.090 1.240 ;
        RECT  12.750 0.840 13.060 2.100 ;
        RECT  12.750 0.450 13.010 2.100 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.058  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.168  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  14.390 1.390 14.550 2.540 ;
        RECT  13.350 1.430 13.510 2.540 ;
        RECT  12.150 1.400 12.350 2.540 ;
        RECT  11.110 1.480 11.310 2.540 ;
        RECT  9.990 2.080 10.270 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  14.330 -0.140 14.610 0.660 ;
        RECT  13.290 -0.140 13.570 0.610 ;
        RECT  12.290 -0.140 12.490 0.610 ;
        RECT  11.270 -0.140 11.430 0.600 ;
        RECT  9.530 -0.140 9.810 0.320 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.100 -0.140 3.300 0.380 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.460 0.720 1.660 1.190 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.620 0.840 ;
        RECT  2.180 0.620 2.400 1.720 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.900 4.960 1.180 ;
        RECT  3.800 0.900 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.820 0.300 2.940 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.780 0.300 2.940 0.700 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  1.820 0.300 2.020 0.680 ;
        RECT  3.460 0.300 3.620 0.700 ;
        RECT  2.780 0.540 3.620 0.700 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.510 0.620 10.790 0.890 ;
        RECT  10.590 1.080 11.610 1.240 ;
        RECT  10.590 0.620 10.790 2.100 ;
        RECT  10.050 0.300 11.110 0.460 ;
        RECT  10.950 0.300 11.110 0.920 ;
        RECT  10.050 0.300 10.210 0.760 ;
        RECT  9.510 0.580 10.090 0.860 ;
        RECT  10.950 0.760 11.970 0.920 ;
        RECT  11.770 0.490 11.970 1.630 ;
        RECT  9.930 0.580 10.090 1.840 ;
        RECT  11.590 1.480 11.950 1.680 ;
        RECT  9.380 1.680 10.090 1.840 ;
        RECT  9.380 1.680 9.660 1.900 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.050 2.400 ;
        RECT  9.970 1.140 14.800 2.400 ;
        RECT  0.000 1.160 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.140 ;
        RECT  9.050 0.000 9.970 1.160 ;
    END
END SDFCQM8HM

MACRO SDFCQM4HM
    CLASS CORE ;
    FOREIGN SDFCQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.060 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.060 3.100 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.591  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.710 0.840 13.110 1.280 ;
        RECT  12.710 0.840 13.030 2.100 ;
        RECT  12.710 0.450 12.970 2.100 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.310 1.400 13.470 2.540 ;
        RECT  12.130 1.410 12.310 2.540 ;
        RECT  11.110 1.480 11.310 2.540 ;
        RECT  9.990 2.080 10.270 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.250 -0.140 13.530 0.660 ;
        RECT  12.250 -0.140 12.450 0.610 ;
        RECT  11.270 -0.140 11.430 0.600 ;
        RECT  9.530 -0.140 9.810 0.320 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.100 -0.140 3.300 0.380 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.460 0.720 1.660 1.190 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.620 0.840 ;
        RECT  2.180 0.620 2.400 1.720 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.940 4.960 1.220 ;
        RECT  3.800 0.940 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.820 0.300 2.940 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.780 0.300 2.940 0.700 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  1.820 0.300 2.020 0.680 ;
        RECT  3.460 0.300 3.620 0.700 ;
        RECT  2.780 0.540 3.620 0.700 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.510 0.620 10.790 0.890 ;
        RECT  10.590 1.080 11.610 1.240 ;
        RECT  10.590 0.620 10.790 2.100 ;
        RECT  10.050 0.300 11.110 0.460 ;
        RECT  10.950 0.300 11.110 0.920 ;
        RECT  10.050 0.300 10.210 0.760 ;
        RECT  9.510 0.580 10.090 0.860 ;
        RECT  10.950 0.760 11.970 0.920 ;
        RECT  11.770 0.490 11.970 1.630 ;
        RECT  9.930 0.580 10.090 1.840 ;
        RECT  11.590 1.480 11.950 1.680 ;
        RECT  9.380 1.680 10.090 1.840 ;
        RECT  9.380 1.680 9.660 1.900 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.010 2.400 ;
        RECT  9.970 1.140 14.000 2.400 ;
        RECT  0.000 1.160 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.140 ;
        RECT  7.010 0.000 9.970 1.160 ;
    END
END SDFCQM4HM

MACRO SDFCQM2HM
    CLASS CORE ;
    FOREIGN SDFCQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.060 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.060 3.100 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.910 0.840 12.300 1.280 ;
        RECT  11.910 0.450 12.110 2.100 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.168  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  12.450 1.420 12.610 2.540 ;
        RECT  10.610 1.480 10.810 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  12.390 -0.140 12.670 0.660 ;
        RECT  10.850 -0.140 11.010 0.600 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.100 -0.140 3.300 0.380 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.460 0.720 1.660 1.190 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.620 0.840 ;
        RECT  2.180 0.620 2.400 1.720 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.940 4.960 1.220 ;
        RECT  3.800 0.940 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.820 0.300 2.940 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.780 0.300 2.940 0.700 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  1.820 0.300 2.020 0.680 ;
        RECT  3.460 0.300 3.620 0.700 ;
        RECT  2.780 0.540 3.620 0.700 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.090 0.620 10.370 1.240 ;
        RECT  10.090 1.080 11.190 1.240 ;
        RECT  10.090 0.620 10.290 2.100 ;
        RECT  9.770 0.300 10.690 0.460 ;
        RECT  10.530 0.300 10.690 0.920 ;
        RECT  9.510 0.580 9.930 0.860 ;
        RECT  10.530 0.760 11.630 0.920 ;
        RECT  11.430 0.300 11.630 1.680 ;
        RECT  11.170 1.480 11.630 1.680 ;
        RECT  9.770 0.300 9.930 1.840 ;
        RECT  9.380 1.680 9.930 1.840 ;
        RECT  9.380 1.680 9.660 1.900 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.010 2.400 ;
        RECT  9.930 1.140 12.800 2.400 ;
        RECT  0.000 1.160 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
        RECT  7.010 0.000 9.930 1.160 ;
    END
END SDFCQM2HM

MACRO SDFCQM1HM
    CLASS CORE ;
    FOREIGN SDFCQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.000 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.120 2.380 1.560 ;
        RECT  1.860 1.120 2.380 1.320 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.910 0.840 12.300 1.280 ;
        RECT  11.910 0.300 12.110 1.720 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.168  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  12.450 1.600 12.610 2.540 ;
        RECT  10.610 1.480 10.810 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  12.390 -0.140 12.670 0.580 ;
        RECT  10.850 -0.140 11.010 0.600 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.020 -0.140 3.300 0.320 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.430 0.800 3.010 0.960 ;
        RECT  1.430 0.720 1.660 1.190 ;
        RECT  2.730 0.800 3.010 1.300 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.940 4.960 1.220 ;
        RECT  3.800 0.940 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.740 0.300 2.860 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.700 0.300 2.860 0.640 ;
        RECT  1.740 0.300 2.100 0.500 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  3.460 0.300 3.620 0.640 ;
        RECT  2.700 0.480 3.620 0.640 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.090 0.620 10.370 1.240 ;
        RECT  10.090 1.080 11.190 1.240 ;
        RECT  10.090 0.620 10.290 2.100 ;
        RECT  9.770 0.300 10.690 0.460 ;
        RECT  10.530 0.300 10.690 0.920 ;
        RECT  9.510 0.580 9.930 0.860 ;
        RECT  10.530 0.760 11.630 0.920 ;
        RECT  11.430 0.300 11.630 1.680 ;
        RECT  11.170 1.480 11.630 1.680 ;
        RECT  9.770 0.300 9.930 1.840 ;
        RECT  9.380 1.680 9.930 1.840 ;
        RECT  9.380 1.680 9.660 1.900 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.010 2.400 ;
        RECT  9.940 1.140 12.800 2.400 ;
        RECT  0.000 1.160 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
        RECT  7.010 0.000 9.940 1.160 ;
    END
END SDFCQM1HM

MACRO SDFCM8HM
    CLASS CORE ;
    FOREIGN SDFCM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.060 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.060 3.100 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.193  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.150 0.460 14.310 1.760 ;
        RECT  12.830 0.840 14.310 1.280 ;
        RECT  12.830 0.450 13.030 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.330 0.380 16.530 2.100 ;
        RECT  15.290 0.840 16.530 1.160 ;
        RECT  15.290 0.380 15.490 2.100 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.058  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.168  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.200 2.540 ;
        RECT  16.850 1.480 17.050 2.540 ;
        RECT  15.810 1.480 16.010 2.540 ;
        RECT  14.790 1.440 14.950 2.540 ;
        RECT  13.510 1.800 13.670 2.540 ;
        RECT  12.150 1.810 12.350 2.540 ;
        RECT  11.110 1.480 11.310 2.540 ;
        RECT  9.990 2.080 10.270 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.200 0.140 ;
        RECT  16.850 -0.140 17.050 0.660 ;
        RECT  15.810 -0.140 16.010 0.660 ;
        RECT  14.670 -0.140 14.950 0.660 ;
        RECT  13.460 -0.140 13.740 0.610 ;
        RECT  12.290 -0.140 12.490 0.610 ;
        RECT  11.270 -0.140 11.430 0.600 ;
        RECT  9.530 -0.140 9.810 0.320 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.100 -0.140 3.300 0.380 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.460 0.720 1.660 1.190 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.620 0.840 ;
        RECT  2.180 0.620 2.400 1.720 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.900 4.960 1.180 ;
        RECT  3.800 0.900 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.820 0.300 2.940 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.780 0.300 2.940 0.700 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  1.820 0.300 2.020 0.680 ;
        RECT  3.460 0.300 3.620 0.700 ;
        RECT  2.780 0.540 3.620 0.700 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.510 0.620 10.790 0.890 ;
        RECT  10.590 1.080 11.610 1.240 ;
        RECT  10.590 0.620 10.790 2.100 ;
        RECT  10.050 0.300 11.110 0.460 ;
        RECT  10.950 0.300 11.110 0.920 ;
        RECT  10.050 0.300 10.210 0.760 ;
        RECT  9.510 0.580 10.090 0.860 ;
        RECT  10.950 0.760 11.970 0.920 ;
        RECT  14.470 1.020 15.030 1.220 ;
        RECT  11.770 0.490 11.970 1.630 ;
        RECT  11.770 1.470 12.670 1.630 ;
        RECT  13.190 1.480 13.990 1.640 ;
        RECT  9.930 0.580 10.090 1.840 ;
        RECT  11.590 1.480 11.950 1.680 ;
        RECT  9.380 1.680 10.090 1.840 ;
        RECT  12.510 1.470 12.670 2.040 ;
        RECT  9.380 1.680 9.660 1.900 ;
        RECT  13.830 1.480 13.990 2.080 ;
        RECT  13.190 1.480 13.350 2.040 ;
        RECT  12.510 1.880 13.350 2.040 ;
        RECT  14.470 1.020 14.630 2.080 ;
        RECT  13.830 1.920 14.630 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.050 2.400 ;
        RECT  9.970 1.140 17.200 2.400 ;
        RECT  0.000 1.160 17.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.200 1.140 ;
        RECT  9.050 0.000 9.970 1.160 ;
    END
END SDFCM8HM

MACRO SDFCM4HM
    CLASS CORE ;
    FOREIGN SDFCM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.060 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.060 3.100 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.616  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.790 0.840 13.110 1.280 ;
        RECT  12.790 0.450 12.990 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.970 0.840 14.400 1.160 ;
        RECT  13.970 0.380 14.170 2.100 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.490 1.480 14.690 2.540 ;
        RECT  13.470 1.800 13.630 2.540 ;
        RECT  12.110 1.810 12.310 2.540 ;
        RECT  11.110 1.480 11.310 2.540 ;
        RECT  9.990 2.080 10.270 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.490 -0.140 14.690 0.660 ;
        RECT  13.350 -0.140 13.630 0.660 ;
        RECT  12.250 -0.140 12.450 0.610 ;
        RECT  11.270 -0.140 11.430 0.600 ;
        RECT  9.530 -0.140 9.810 0.320 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.100 -0.140 3.300 0.380 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.460 0.720 1.660 1.190 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.620 0.840 ;
        RECT  2.180 0.620 2.400 1.720 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.940 4.960 1.220 ;
        RECT  3.800 0.940 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.820 0.300 2.940 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.780 0.300 2.940 0.700 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  1.820 0.300 2.020 0.680 ;
        RECT  3.460 0.300 3.620 0.700 ;
        RECT  2.780 0.540 3.620 0.700 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.510 0.620 10.790 0.890 ;
        RECT  10.590 1.080 11.610 1.240 ;
        RECT  10.590 0.620 10.790 2.100 ;
        RECT  10.050 0.300 11.110 0.460 ;
        RECT  10.950 0.300 11.110 0.920 ;
        RECT  10.050 0.300 10.210 0.760 ;
        RECT  9.510 0.580 10.090 0.860 ;
        RECT  10.950 0.760 11.970 0.920 ;
        RECT  13.370 1.020 13.710 1.220 ;
        RECT  11.770 0.490 11.970 1.630 ;
        RECT  11.770 1.470 12.630 1.630 ;
        RECT  13.370 1.020 13.530 1.640 ;
        RECT  13.150 1.480 13.530 1.640 ;
        RECT  9.930 0.580 10.090 1.840 ;
        RECT  11.590 1.480 11.950 1.680 ;
        RECT  9.380 1.680 10.090 1.840 ;
        RECT  12.470 1.470 12.630 2.040 ;
        RECT  9.380 1.680 9.660 1.900 ;
        RECT  13.150 1.480 13.310 2.040 ;
        RECT  12.470 1.880 13.310 2.040 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.010 2.400 ;
        RECT  9.970 1.140 15.200 2.400 ;
        RECT  0.000 1.160 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 1.140 ;
        RECT  7.010 0.000 9.970 1.160 ;
    END
END SDFCM4HM

MACRO SDFCM2HM
    CLASS CORE ;
    FOREIGN SDFCM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.060 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.060 3.100 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.910 0.840 12.300 1.280 ;
        RECT  11.910 0.450 12.110 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.090 0.840 13.500 1.160 ;
        RECT  13.090 0.380 13.290 2.100 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.168  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.590 1.800 12.750 2.540 ;
        RECT  10.610 1.480 10.810 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.470 -0.140 12.750 0.660 ;
        RECT  10.850 -0.140 11.010 0.600 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.100 -0.140 3.300 0.380 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.460 0.720 1.660 1.190 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.180 0.620 2.620 0.840 ;
        RECT  2.180 0.620 2.400 1.720 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.940 4.960 1.220 ;
        RECT  3.800 0.940 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.820 0.300 2.940 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.780 0.300 2.940 0.700 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  1.820 0.300 2.020 0.680 ;
        RECT  3.460 0.300 3.620 0.700 ;
        RECT  2.780 0.540 3.620 0.700 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.090 0.620 10.370 1.240 ;
        RECT  10.090 1.080 11.190 1.240 ;
        RECT  10.090 0.620 10.290 2.100 ;
        RECT  9.770 0.300 10.690 0.460 ;
        RECT  10.530 0.300 10.690 0.920 ;
        RECT  9.510 0.580 9.930 0.860 ;
        RECT  10.530 0.760 11.630 0.920 ;
        RECT  12.770 0.940 12.930 1.640 ;
        RECT  12.270 1.480 12.930 1.640 ;
        RECT  11.170 1.480 11.630 1.680 ;
        RECT  9.770 0.300 9.930 1.840 ;
        RECT  9.380 1.680 9.930 1.840 ;
        RECT  11.430 0.300 11.630 2.040 ;
        RECT  11.390 1.480 11.630 2.040 ;
        RECT  9.380 1.680 9.660 1.900 ;
        RECT  12.270 1.480 12.430 2.040 ;
        RECT  11.390 1.880 12.430 2.040 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.010 2.400 ;
        RECT  9.930 1.140 13.600 2.400 ;
        RECT  0.000 1.160 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.140 ;
        RECT  7.010 0.000 9.930 1.160 ;
    END
END SDFCM2HM

MACRO SDFCM1HM
    CLASS CORE ;
    FOREIGN SDFCM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.000 3.610 1.560 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.120 2.380 1.560 ;
        RECT  1.860 1.120 2.380 1.320 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.910 0.840 12.300 1.280 ;
        RECT  11.910 0.300 12.110 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.090 0.840 13.500 1.160 ;
        RECT  13.090 0.300 13.290 2.010 ;
        END
    END QB
    PIN SD
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.180 1.560 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.168  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.590 1.800 12.750 2.540 ;
        RECT  10.610 1.480 10.810 2.540 ;
        RECT  7.380 1.760 7.580 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.470 -0.140 12.750 0.580 ;
        RECT  10.850 -0.140 11.010 0.600 ;
        RECT  7.150 -0.140 7.430 0.320 ;
        RECT  4.560 -0.140 4.760 0.420 ;
        RECT  3.020 -0.140 3.300 0.320 ;
        RECT  0.700 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 1.660 0.880 ;
        RECT  1.430 0.800 3.010 0.960 ;
        RECT  1.430 0.720 1.660 1.190 ;
        RECT  2.730 0.800 3.010 1.300 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  3.800 0.620 4.080 1.660 ;
        RECT  3.800 0.940 4.960 1.220 ;
        RECT  3.800 0.940 4.120 1.660 ;
        RECT  1.680 1.480 1.880 2.040 ;
        RECT  2.560 1.760 3.600 1.920 ;
        RECT  1.680 1.880 2.720 2.040 ;
        RECT  3.440 1.840 5.750 2.040 ;
        RECT  1.740 0.300 2.860 0.460 ;
        RECT  3.460 0.300 4.400 0.460 ;
        RECT  4.920 0.300 5.970 0.460 ;
        RECT  2.700 0.300 2.860 0.640 ;
        RECT  1.740 0.300 2.100 0.500 ;
        RECT  4.240 0.300 4.400 0.740 ;
        RECT  3.460 0.300 3.620 0.640 ;
        RECT  2.700 0.480 3.620 0.640 ;
        RECT  4.920 0.300 5.080 0.740 ;
        RECT  4.240 0.580 5.080 0.740 ;
        RECT  5.770 0.300 5.970 0.780 ;
        RECT  5.240 0.620 5.520 1.660 ;
        RECT  4.740 1.500 6.070 1.660 ;
        RECT  5.910 1.500 6.070 2.100 ;
        RECT  5.910 1.940 6.980 2.100 ;
        RECT  6.250 0.420 6.480 1.780 ;
        RECT  6.230 1.120 6.480 1.780 ;
        RECT  7.600 1.120 7.800 1.520 ;
        RECT  6.230 1.360 7.800 1.520 ;
        RECT  6.230 1.360 6.510 1.780 ;
        RECT  7.940 0.620 8.220 0.960 ;
        RECT  7.120 0.800 8.220 0.960 ;
        RECT  7.120 0.800 7.320 1.200 ;
        RECT  7.960 0.620 8.160 1.890 ;
        RECT  8.620 0.620 8.980 0.840 ;
        RECT  8.620 0.620 8.900 1.810 ;
        RECT  8.680 1.640 8.960 2.100 ;
        RECT  7.590 0.300 9.310 0.460 ;
        RECT  6.640 0.300 6.920 0.640 ;
        RECT  7.590 0.300 7.750 0.640 ;
        RECT  6.640 0.480 7.750 0.640 ;
        RECT  9.140 0.300 9.310 1.460 ;
        RECT  9.140 1.240 9.610 1.460 ;
        RECT  10.090 0.620 10.370 1.240 ;
        RECT  10.090 1.080 11.190 1.240 ;
        RECT  10.090 0.620 10.290 2.100 ;
        RECT  9.770 0.300 10.690 0.460 ;
        RECT  10.530 0.300 10.690 0.920 ;
        RECT  9.510 0.580 9.930 0.860 ;
        RECT  10.530 0.760 11.630 0.920 ;
        RECT  12.770 0.940 12.930 1.640 ;
        RECT  12.270 1.480 12.930 1.640 ;
        RECT  11.170 1.480 11.630 1.680 ;
        RECT  9.770 0.300 9.930 1.840 ;
        RECT  9.380 1.680 9.930 1.840 ;
        RECT  11.430 0.300 11.630 2.040 ;
        RECT  11.390 1.480 11.630 2.040 ;
        RECT  9.380 1.680 9.660 1.900 ;
        RECT  12.270 1.480 12.430 2.040 ;
        RECT  11.390 1.880 12.430 2.040 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.010 2.400 ;
        RECT  9.940 1.140 13.600 2.400 ;
        RECT  0.000 1.160 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.140 ;
        RECT  7.010 0.000 9.940 1.160 ;
    END
END SDFCM1HM

MACRO OR6M8HM
    CLASS CORE ;
    FOREIGN OR6M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.347  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.610 1.480 8.810 1.960 ;
        RECT  4.450 1.480 8.810 1.680 ;
        RECT  6.900 0.700 8.330 0.880 ;
        RECT  8.050 0.660 8.330 0.880 ;
        RECT  7.570 1.480 7.770 1.960 ;
        RECT  6.900 0.660 7.290 0.880 ;
        RECT  6.900 0.660 7.100 1.680 ;
        RECT  6.530 1.480 6.730 1.960 ;
        RECT  5.490 1.480 5.690 1.960 ;
        RECT  4.450 1.480 4.650 1.960 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.602  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.700 1.000 9.900 1.200 ;
        LAYER ME2 ;
        RECT  9.700 0.800 9.900 1.350 ;
        LAYER ME1 ;
        RECT  9.450 1.000 10.030 1.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.828  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  11.300 1.000 11.500 1.200 ;
        LAYER ME2 ;
        RECT  11.300 0.800 11.500 1.350 ;
        LAYER ME1 ;
        RECT  10.910 1.000 11.600 1.200 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.725  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  12.100 1.000 12.300 1.200 ;
        LAYER ME2 ;
        RECT  12.100 0.800 12.300 1.350 ;
        LAYER ME1 ;
        RECT  11.950 1.000 12.590 1.200 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.664  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.000 3.500 1.200 ;
        LAYER ME2 ;
        RECT  3.300 0.800 3.500 1.350 ;
        LAYER ME1 ;
        RECT  3.200 1.000 3.810 1.200 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.828  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.000 2.300 1.200 ;
        LAYER ME2 ;
        RECT  2.100 0.800 2.300 1.350 ;
        LAYER ME1 ;
        RECT  1.710 1.000 2.400 1.200 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.725  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.000 1.100 1.200 ;
        LAYER ME2 ;
        RECT  0.900 0.800 1.100 1.350 ;
        LAYER ME1 ;
        RECT  0.670 1.000 1.310 1.200 ;
        END
    END F
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.170 1.800 12.370 2.540 ;
        RECT  8.090 1.840 8.290 2.540 ;
        RECT  7.050 1.840 7.250 2.540 ;
        RECT  6.010 1.840 6.210 2.540 ;
        RECT  4.970 1.840 5.170 2.540 ;
        RECT  0.890 1.840 1.090 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.690 -0.140 12.890 0.570 ;
        RECT  11.610 -0.140 11.890 0.500 ;
        RECT  10.570 -0.140 10.850 0.500 ;
        RECT  10.090 -0.140 10.370 0.500 ;
        RECT  9.050 -0.140 9.330 0.500 ;
        RECT  6.010 -0.140 6.210 0.600 ;
        RECT  4.970 -0.140 5.170 0.600 ;
        RECT  3.930 -0.140 4.210 0.500 ;
        RECT  2.890 -0.140 3.170 0.500 ;
        RECT  2.410 -0.140 2.690 0.500 ;
        RECT  1.370 -0.140 1.650 0.500 ;
        RECT  0.370 -0.140 0.570 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.370 1.440 2.690 1.640 ;
        RECT  0.370 1.440 0.570 2.080 ;
        RECT  1.410 1.440 1.610 2.080 ;
        RECT  1.890 1.880 3.690 2.080 ;
        RECT  0.890 0.320 1.090 0.820 ;
        RECT  1.930 0.320 2.130 0.820 ;
        RECT  3.450 0.300 3.650 0.820 ;
        RECT  0.890 0.660 4.170 0.820 ;
        RECT  3.970 1.100 6.110 1.300 ;
        RECT  2.890 1.500 4.170 1.700 ;
        RECT  3.970 0.660 4.170 2.080 ;
        RECT  6.530 0.340 8.810 0.500 ;
        RECT  7.530 0.340 7.810 0.540 ;
        RECT  8.610 0.340 8.810 0.620 ;
        RECT  4.450 0.380 4.650 0.920 ;
        RECT  5.490 0.470 5.690 0.920 ;
        RECT  6.530 0.340 6.730 0.920 ;
        RECT  4.450 0.760 6.730 0.920 ;
        RECT  9.570 1.880 11.370 2.080 ;
        RECT  9.610 0.300 9.810 0.830 ;
        RECT  11.130 0.320 11.330 0.830 ;
        RECT  12.170 0.320 12.370 0.830 ;
        RECT  9.090 0.660 12.370 0.830 ;
        RECT  7.460 1.100 9.290 1.300 ;
        RECT  9.090 1.520 10.370 1.720 ;
        RECT  9.090 0.660 9.290 2.080 ;
        RECT  10.570 1.440 12.890 1.640 ;
        RECT  11.650 1.440 11.850 2.080 ;
        RECT  12.690 1.440 12.890 2.080 ;
        LAYER VTPH ;
        RECT  8.940 1.100 13.200 2.400 ;
        RECT  0.000 1.100 4.280 2.400 ;
        RECT  8.940 1.140 13.600 2.400 ;
        RECT  0.000 1.180 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.100 ;
        RECT  13.200 0.000 13.600 1.140 ;
        RECT  4.280 0.000 8.940 1.180 ;
    END
END OR6M8HM

MACRO OR6M6HM
    CLASS CORE ;
    FOREIGN OR6M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.212  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.922  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.040 1.000 3.240 1.200 ;
        RECT  1.400 1.000 1.600 1.200 ;
        LAYER ME2 ;
        RECT  3.040 0.540 3.240 1.260 ;
        RECT  1.400 0.540 3.240 0.740 ;
        RECT  1.300 0.840 1.600 1.310 ;
        RECT  1.400 0.540 1.600 1.310 ;
        LAYER ME1 ;
        RECT  2.980 1.000 3.600 1.200 ;
        RECT  1.100 1.000 1.790 1.200 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        ANTENNAGATEAREA 0.212  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.827  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.620 1.080 9.820 1.280 ;
        LAYER ME2 ;
        RECT  9.620 0.840 9.900 1.380 ;
        LAYER ME1 ;
        RECT  7.740 1.080 9.920 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        ANTENNAGATEAREA 0.212  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.959  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.300 0.720 8.500 0.920 ;
        LAYER ME2 ;
        RECT  8.100 0.620 8.500 1.160 ;
        LAYER ME1 ;
        RECT  8.000 0.720 8.600 0.920 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.720 0.840 11.100 1.300 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.900 0.320 1.630 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.998  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.840 0.740 7.140 0.900 ;
        RECT  6.980 0.400 7.140 0.900 ;
        RECT  6.440 1.480 6.640 2.020 ;
        RECT  4.360 1.480 6.640 1.680 ;
        RECT  5.840 0.740 6.300 1.680 ;
        RECT  5.840 0.620 6.200 1.680 ;
        RECT  5.400 1.480 5.600 2.020 ;
        RECT  4.360 1.480 4.560 2.060 ;
        END
    END Z
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        ANTENNAGATEAREA 0.212  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.326  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.000 2.300 1.200 ;
        LAYER ME2 ;
        RECT  2.100 0.940 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.990 1.000 2.740 1.200 ;
        END
    END F
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  8.680 2.080 8.960 2.540 ;
        RECT  6.960 1.740 7.160 2.540 ;
        RECT  5.920 1.840 6.120 2.540 ;
        RECT  4.880 1.840 5.080 2.540 ;
        RECT  3.840 1.780 4.040 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.500 -0.140 10.780 0.500 ;
        RECT  9.340 -0.140 9.620 0.500 ;
        RECT  4.840 -0.140 5.120 0.500 ;
        RECT  3.800 -0.140 4.080 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.660 1.700 3.080 1.900 ;
        RECT  1.180 1.360 3.560 1.520 ;
        RECT  0.140 1.820 0.340 2.100 ;
        RECT  3.360 1.360 3.560 1.960 ;
        RECT  1.180 1.360 1.380 2.100 ;
        RECT  0.140 1.940 1.380 2.100 ;
        RECT  1.180 0.430 1.380 0.820 ;
        RECT  2.220 0.450 2.420 0.820 ;
        RECT  0.490 0.660 4.000 0.820 ;
        RECT  3.840 0.660 4.000 1.220 ;
        RECT  3.840 1.020 5.140 1.220 ;
        RECT  0.490 0.660 0.650 1.760 ;
        RECT  0.490 1.560 0.900 1.760 ;
        RECT  5.400 0.300 6.640 0.460 ;
        RECT  6.440 0.300 6.640 0.580 ;
        RECT  4.360 0.380 4.560 0.860 ;
        RECT  5.400 0.300 5.600 0.860 ;
        RECT  4.360 0.660 5.600 0.860 ;
        RECT  7.920 1.440 9.740 1.600 ;
        RECT  7.920 1.440 8.200 1.740 ;
        RECT  9.460 1.440 9.740 1.740 ;
        RECT  7.300 0.300 8.960 0.460 ;
        RECT  8.760 0.300 8.960 0.820 ;
        RECT  10.020 0.430 10.220 0.820 ;
        RECT  8.760 0.660 10.460 0.820 ;
        RECT  7.300 0.300 7.460 1.310 ;
        RECT  6.580 1.110 7.460 1.310 ;
        RECT  10.260 0.660 10.460 1.740 ;
        RECT  10.260 1.580 10.820 1.740 ;
        RECT  8.360 1.760 9.300 1.920 ;
        RECT  7.360 1.900 8.520 2.060 ;
        RECT  11.060 1.690 11.260 2.060 ;
        RECT  9.120 1.900 11.260 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.140 ;
    END
END OR6M6HM

MACRO OR6M4HM
    CLASS CORE ;
    FOREIGN OR6M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        ANTENNAGATEAREA 0.122  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.399  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.850 1.000 5.050 1.200 ;
        LAYER ME2 ;
        RECT  4.850 0.840 5.100 1.300 ;
        LAYER ME1 ;
        RECT  4.650 1.000 5.250 1.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.570 1.080 5.900 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 1.040 6.330 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.990 1.550 1.560 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.040 1.100 1.560 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.160 ;
        END
    END F
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.616  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.620 3.990 2.010 ;
        RECT  2.710 1.580 3.990 1.740 ;
        RECT  2.710 1.580 2.910 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.310 1.840 6.510 2.540 ;
        RECT  4.230 1.900 4.510 2.540 ;
        RECT  3.190 1.900 3.470 2.540 ;
        RECT  2.190 1.740 2.390 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.310 -0.140 6.510 0.590 ;
        RECT  5.230 -0.140 5.510 0.500 ;
        RECT  2.670 -0.140 2.950 0.500 ;
        RECT  1.150 -0.140 1.430 0.500 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.310 0.860 0.820 ;
        RECT  0.660 0.660 1.910 0.820 ;
        RECT  1.710 1.080 3.130 1.280 ;
        RECT  1.710 0.310 1.910 2.100 ;
        RECT  3.230 0.300 4.510 0.460 ;
        RECT  4.230 0.300 4.510 0.520 ;
        RECT  2.190 0.420 2.390 0.860 ;
        RECT  3.230 0.300 3.430 0.860 ;
        RECT  2.190 0.660 3.430 0.860 ;
        RECT  4.750 0.310 4.950 0.840 ;
        RECT  5.790 0.310 5.990 0.840 ;
        RECT  4.150 0.680 5.990 0.840 ;
        RECT  4.150 0.680 4.350 1.740 ;
        RECT  4.150 1.540 4.950 1.740 ;
        RECT  4.750 1.540 4.950 1.970 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END OR6M4HM

MACRO OR6M2HM
    CLASS CORE ;
    FOREIGN OR6M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.810 1.050 1.010 1.250 ;
        LAYER ME2 ;
        RECT  0.810 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.730 0.950 1.050 1.350 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.634  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.120 1.130 4.320 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.320 1.430 ;
        LAYER ME1 ;
        RECT  4.120 1.000 4.440 1.450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.815  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.640 1.000 3.840 1.200 ;
        LAYER ME2 ;
        RECT  3.580 0.840 3.900 1.310 ;
        LAYER ME1 ;
        RECT  3.470 1.000 3.960 1.310 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.700 1.160 5.100 1.620 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 0.900 1.960 1.100 ;
        RECT  1.560 0.900 1.840 1.200 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.400 1.560 ;
        END
    END F
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.386  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.320 3.100 0.520 ;
        RECT  2.500 1.860 2.780 2.060 ;
        RECT  2.500 0.320 2.700 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.700 1.840 4.900 2.540 ;
        RECT  3.020 1.900 3.300 2.540 ;
        RECT  1.980 1.840 2.200 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.860 -0.140 5.060 0.840 ;
        RECT  3.860 -0.140 4.060 0.840 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.540 0.720 ;
        RECT  1.210 0.520 1.370 2.050 ;
        RECT  2.040 1.310 2.320 1.680 ;
        RECT  1.210 1.520 2.320 1.680 ;
        RECT  1.210 1.520 1.550 2.050 ;
        RECT  3.300 0.560 3.580 0.840 ;
        RECT  2.900 0.680 3.580 0.840 ;
        RECT  2.900 0.680 3.100 1.740 ;
        RECT  2.900 1.540 3.740 1.740 ;
        RECT  3.540 1.540 3.740 1.970 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OR6M2HM

MACRO OR6M1HM
    CLASS CORE ;
    FOREIGN OR6M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.815  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.640 1.000 3.840 1.200 ;
        LAYER ME2 ;
        RECT  3.580 0.840 3.900 1.310 ;
        LAYER ME1 ;
        RECT  3.470 1.000 3.960 1.310 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.634  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.120 1.130 4.320 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.320 1.430 ;
        LAYER ME1 ;
        RECT  4.120 1.000 4.440 1.450 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.810 1.050 1.010 1.250 ;
        LAYER ME2 ;
        RECT  0.810 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.730 0.950 1.050 1.350 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.700 1.160 5.100 1.620 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 0.900 1.960 1.100 ;
        RECT  1.560 0.900 1.840 1.200 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.400 1.560 ;
        END
    END F
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.269  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.320 3.100 0.520 ;
        RECT  2.500 1.860 2.780 2.060 ;
        RECT  2.500 0.320 2.700 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.700 1.840 4.900 2.540 ;
        RECT  3.020 1.900 3.300 2.540 ;
        RECT  1.980 1.840 2.200 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.860 -0.140 5.060 0.840 ;
        RECT  3.860 -0.140 4.060 0.840 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.540 0.720 ;
        RECT  1.210 0.520 1.370 2.050 ;
        RECT  2.040 1.310 2.320 1.680 ;
        RECT  1.210 1.520 2.320 1.680 ;
        RECT  1.210 1.520 1.550 2.050 ;
        RECT  3.300 0.560 3.580 0.840 ;
        RECT  2.900 0.680 3.580 0.840 ;
        RECT  2.900 0.680 3.100 1.740 ;
        RECT  2.900 1.540 3.740 1.740 ;
        RECT  3.540 1.540 3.740 1.970 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OR6M1HM

MACRO OR6M12HM
    CLASS CORE ;
    FOREIGN OR6M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  12.100 1.000 12.300 1.200 ;
        LAYER ME2 ;
        RECT  12.100 0.800 12.300 1.350 ;
        LAYER ME1 ;
        RECT  11.700 1.000 12.700 1.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  13.300 1.000 13.500 1.200 ;
        LAYER ME2 ;
        RECT  13.300 0.800 13.500 1.350 ;
        LAYER ME1 ;
        RECT  13.100 1.000 14.100 1.200 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.860  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.640 0.660 10.960 0.860 ;
        RECT  10.760 0.430 10.960 0.860 ;
        RECT  10.240 1.480 10.440 1.960 ;
        RECT  6.080 1.480 10.440 1.680 ;
        RECT  9.200 1.480 9.400 1.960 ;
        RECT  8.640 0.660 9.100 1.680 ;
        RECT  8.160 1.480 8.360 1.960 ;
        RECT  7.120 1.480 7.320 1.960 ;
        RECT  6.080 1.480 6.280 1.960 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  14.900 1.000 15.100 1.200 ;
        LAYER ME2 ;
        RECT  14.900 0.800 15.100 1.350 ;
        LAYER ME1 ;
        RECT  14.660 1.000 15.660 1.200 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.000 4.300 1.200 ;
        LAYER ME2 ;
        RECT  4.100 0.800 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.820 1.000 4.820 1.200 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.000 2.700 1.200 ;
        LAYER ME2 ;
        RECT  2.500 0.800 2.700 1.350 ;
        LAYER ME1 ;
        RECT  2.260 1.000 3.260 1.200 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.000 1.100 1.200 ;
        LAYER ME2 ;
        RECT  0.900 0.800 1.100 1.350 ;
        LAYER ME1 ;
        RECT  0.700 1.000 1.700 1.200 ;
        END
    END F
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.800 2.540 ;
        RECT  15.920 1.440 16.120 2.540 ;
        RECT  14.880 1.800 15.080 2.540 ;
        RECT  10.760 1.680 10.960 2.540 ;
        RECT  9.720 1.840 9.920 2.540 ;
        RECT  8.680 1.840 8.880 2.540 ;
        RECT  7.640 1.840 7.840 2.540 ;
        RECT  6.600 1.840 6.800 2.540 ;
        RECT  5.560 1.680 5.760 2.540 ;
        RECT  1.440 1.840 1.640 2.540 ;
        RECT  0.400 1.480 0.600 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.800 0.140 ;
        RECT  15.400 -0.140 15.600 0.640 ;
        RECT  14.320 -0.140 14.600 0.500 ;
        RECT  13.280 -0.140 13.560 0.500 ;
        RECT  12.240 -0.140 12.520 0.500 ;
        RECT  11.200 -0.140 11.480 0.500 ;
        RECT  7.640 -0.140 7.840 0.560 ;
        RECT  6.600 -0.140 6.800 0.560 ;
        RECT  5.560 -0.140 5.760 0.710 ;
        RECT  5.040 -0.140 5.320 0.500 ;
        RECT  4.000 -0.140 4.280 0.500 ;
        RECT  2.960 -0.140 3.240 0.500 ;
        RECT  1.920 -0.140 2.200 0.500 ;
        RECT  0.920 -0.140 1.120 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.920 1.440 3.240 1.640 ;
        RECT  0.920 1.440 1.120 2.080 ;
        RECT  1.960 1.440 2.160 2.080 ;
        RECT  3.520 1.440 3.720 2.080 ;
        RECT  3.520 1.860 4.800 2.080 ;
        RECT  2.440 1.880 4.800 2.080 ;
        RECT  1.440 0.360 1.640 0.820 ;
        RECT  2.480 0.360 2.680 0.820 ;
        RECT  4.560 0.360 4.760 0.820 ;
        RECT  1.440 0.660 5.280 0.820 ;
        RECT  5.080 1.100 7.940 1.300 ;
        RECT  4.000 1.500 5.280 1.700 ;
        RECT  5.080 0.660 5.280 2.080 ;
        RECT  8.160 0.340 10.520 0.500 ;
        RECT  6.080 0.430 6.280 0.920 ;
        RECT  7.120 0.430 7.320 0.920 ;
        RECT  8.160 0.340 8.360 0.920 ;
        RECT  6.080 0.720 8.360 0.920 ;
        RECT  12.800 1.440 13.000 2.080 ;
        RECT  11.720 1.880 14.080 2.080 ;
        RECT  11.760 0.430 11.960 0.830 ;
        RECT  13.840 0.430 14.040 0.830 ;
        RECT  14.880 0.430 15.080 0.830 ;
        RECT  11.240 0.660 15.080 0.830 ;
        RECT  9.520 1.100 11.440 1.300 ;
        RECT  11.240 1.520 12.520 1.720 ;
        RECT  11.240 0.660 11.440 2.080 ;
        RECT  13.280 1.440 15.600 1.640 ;
        RECT  14.360 1.440 14.560 2.080 ;
        RECT  15.400 1.440 15.600 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.080 5.410 2.400 ;
        RECT  11.090 1.080 16.800 2.400 ;
        RECT  0.000 1.180 16.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.800 1.080 ;
        RECT  5.410 0.000 11.090 1.180 ;
    END
END OR6M12HM

MACRO OR6M0HM
    CLASS CORE ;
    FOREIGN OR6M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.810 1.050 1.010 1.250 ;
        LAYER ME2 ;
        RECT  0.810 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.730 0.950 1.050 1.350 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.634  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.120 1.130 4.320 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.320 1.430 ;
        LAYER ME1 ;
        RECT  4.120 1.000 4.440 1.450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.815  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.640 1.000 3.840 1.200 ;
        LAYER ME2 ;
        RECT  3.580 0.840 3.900 1.310 ;
        LAYER ME1 ;
        RECT  3.470 1.000 3.960 1.310 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.700 1.160 5.100 1.620 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 0.900 1.960 1.100 ;
        RECT  1.560 0.900 1.840 1.200 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.400 1.560 ;
        END
    END F
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.217  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.320 3.100 0.520 ;
        RECT  2.500 1.880 2.780 2.080 ;
        RECT  2.500 0.320 2.700 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.700 1.840 4.900 2.540 ;
        RECT  3.020 1.900 3.300 2.540 ;
        RECT  1.980 1.840 2.200 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.860 -0.140 5.060 0.840 ;
        RECT  3.860 -0.140 4.060 0.840 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.540 0.720 ;
        RECT  1.210 0.520 1.370 2.050 ;
        RECT  2.040 1.310 2.320 1.680 ;
        RECT  1.210 1.520 2.320 1.680 ;
        RECT  1.210 1.520 1.550 2.050 ;
        RECT  3.300 0.560 3.580 0.840 ;
        RECT  2.900 0.680 3.580 0.840 ;
        RECT  2.900 0.680 3.100 1.740 ;
        RECT  2.900 1.540 3.740 1.740 ;
        RECT  3.540 1.540 3.740 1.970 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OR6M0HM

MACRO OR4M8HM
    CLASS CORE ;
    FOREIGN OR4M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.076  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.870 1.120 3.070 1.320 ;
        LAYER ME2 ;
        RECT  2.850 0.840 3.100 1.450 ;
        LAYER ME1 ;
        RECT  2.520 1.120 3.240 1.320 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.076  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.000 1.120 1.200 1.320 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.220 1.450 ;
        LAYER ME1 ;
        RECT  0.720 1.120 1.440 1.320 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.440 0.800 3.640 1.260 ;
        RECT  2.100 0.800 3.640 0.960 ;
        RECT  2.100 0.800 2.320 1.260 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.800 1.840 1.260 ;
        RECT  0.100 0.800 1.840 0.960 ;
        RECT  0.100 0.800 0.520 1.300 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.660 0.350 5.900 2.080 ;
        RECT  4.620 1.440 5.900 1.640 ;
        RECT  4.620 0.660 5.900 0.860 ;
        RECT  4.620 1.440 4.820 2.080 ;
        RECT  4.620 0.390 4.820 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.180 1.480 6.380 2.540 ;
        RECT  5.100 1.900 5.380 2.540 ;
        RECT  4.120 1.440 4.280 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.180 -0.140 6.380 0.670 ;
        RECT  5.100 -0.140 5.380 0.500 ;
        RECT  4.120 -0.140 4.280 0.700 ;
        RECT  2.940 -0.140 3.220 0.320 ;
        RECT  1.820 -0.140 2.100 0.320 ;
        RECT  0.780 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.500 2.070 1.700 ;
        RECT  1.870 1.500 2.070 2.080 ;
        RECT  1.870 1.880 3.860 2.080 ;
        RECT  1.220 0.480 3.960 0.640 ;
        RECT  3.800 1.040 5.400 1.240 ;
        RECT  3.800 0.480 3.960 1.720 ;
        RECT  2.700 1.560 3.960 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END OR4M8HM

MACRO OR4M6HM
    CLASS CORE ;
    FOREIGN OR4M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.076  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.780 1.120 2.980 1.320 ;
        LAYER ME2 ;
        RECT  2.780 0.840 3.160 1.450 ;
        LAYER ME1 ;
        RECT  2.520 1.120 3.240 1.320 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.076  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.000 1.120 1.200 1.320 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.220 1.450 ;
        LAYER ME1 ;
        RECT  0.720 1.120 1.440 1.320 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.440 0.800 3.640 1.260 ;
        RECT  2.100 0.800 3.640 0.960 ;
        RECT  2.100 0.800 2.320 1.260 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.800 1.840 1.260 ;
        RECT  0.100 0.800 1.840 0.960 ;
        RECT  0.100 0.800 0.520 1.300 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.660 0.350 5.900 2.080 ;
        RECT  4.620 1.440 5.900 1.640 ;
        RECT  4.620 0.660 5.900 0.860 ;
        RECT  4.620 1.440 4.820 2.080 ;
        RECT  4.620 0.390 4.820 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.100 1.900 5.380 2.540 ;
        RECT  4.120 1.440 4.280 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.380 0.500 ;
        RECT  4.120 -0.140 4.280 0.700 ;
        RECT  2.940 -0.140 3.220 0.320 ;
        RECT  1.820 -0.140 2.100 0.320 ;
        RECT  0.780 -0.140 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.500 2.070 1.700 ;
        RECT  1.870 1.500 2.070 2.080 ;
        RECT  1.870 1.880 3.860 2.080 ;
        RECT  1.220 0.480 3.960 0.640 ;
        RECT  3.800 1.040 5.400 1.240 ;
        RECT  3.800 0.480 3.960 1.720 ;
        RECT  2.700 1.560 3.960 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END OR4M6HM

MACRO OR4M4HM
    CLASS CORE ;
    FOREIGN OR4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 1.060 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.120 1.400 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.020 1.700 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.116  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.960 0.840 2.300 1.220 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.060 1.460 3.500 1.660 ;
        RECT  3.300 0.660 3.500 1.660 ;
        RECT  3.060 0.660 3.500 0.860 ;
        RECT  3.060 1.460 3.260 2.100 ;
        RECT  3.060 0.350 3.260 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.540 1.900 3.820 2.540 ;
        RECT  2.540 1.810 2.740 2.540 ;
        RECT  2.200 1.800 2.360 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.540 -0.140 3.820 0.500 ;
        RECT  2.460 -0.140 2.740 0.320 ;
        RECT  1.260 -0.140 1.540 0.320 ;
        RECT  0.140 -0.140 0.340 0.830 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.520 2.620 0.680 ;
        RECT  2.460 1.020 3.120 1.220 ;
        RECT  2.460 0.520 2.620 1.640 ;
        RECT  1.860 1.480 2.620 1.640 ;
        RECT  1.860 1.480 2.020 2.010 ;
        RECT  0.100 1.810 2.020 2.010 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END OR4M4HM

MACRO OR4M2HM
    CLASS CORE ;
    FOREIGN OR4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.100 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.080 1.100 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.080 1.680 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.880 1.080 2.300 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 0.350 3.100 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.100 2.080 2.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.300 -0.140 2.580 0.500 ;
        RECT  1.180 -0.140 1.460 0.540 ;
        RECT  0.140 -0.140 0.340 0.840 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.610 0.620 0.900 0.920 ;
        RECT  1.740 0.620 2.020 0.920 ;
        RECT  0.610 0.760 2.640 0.920 ;
        RECT  2.460 0.760 2.640 1.920 ;
        RECT  0.100 1.720 2.640 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OR4M2HM

MACRO OR4M1HM
    CLASS CORE ;
    FOREIGN OR4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.100 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.080 1.100 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.080 1.680 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.880 1.080 2.300 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 0.340 3.100 1.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.100 2.080 2.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.300 -0.140 2.580 0.540 ;
        RECT  1.180 -0.140 1.460 0.540 ;
        RECT  0.140 -0.140 0.340 0.840 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.610 0.620 0.900 0.920 ;
        RECT  1.740 0.620 2.020 0.920 ;
        RECT  0.610 0.760 2.640 0.920 ;
        RECT  2.460 0.760 2.640 1.920 ;
        RECT  0.100 1.720 2.640 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OR4M1HM

MACRO OR4M16HM
    CLASS CORE ;
    FOREIGN OR4M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.372  LAYER ME1  ;
        ANTENNAGATEAREA 0.372  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.020 2.700 1.220 ;
        LAYER ME2 ;
        RECT  2.500 0.800 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.000 1.020 3.000 1.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.372  LAYER ME1  ;
        ANTENNAGATEAREA 0.372  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.800 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.500 1.020 1.500 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.888  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.020 1.440 10.220 2.080 ;
        RECT  6.900 0.660 10.220 0.860 ;
        RECT  10.020 0.380 10.220 0.860 ;
        RECT  6.900 1.440 10.220 1.630 ;
        RECT  8.980 1.440 9.180 2.080 ;
        RECT  8.980 0.380 9.180 0.860 ;
        RECT  6.900 1.440 9.180 1.640 ;
        RECT  8.450 0.660 8.750 1.640 ;
        RECT  7.940 1.440 8.140 2.080 ;
        RECT  7.940 0.380 8.140 0.860 ;
        RECT  6.900 1.440 7.100 2.080 ;
        RECT  6.900 0.380 7.100 0.860 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.372  LAYER ME1  ;
        ANTENNAGATEAREA 0.372  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.020 3.900 1.220 ;
        LAYER ME2 ;
        RECT  3.700 0.800 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.560 1.020 4.560 1.220 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.372  LAYER ME1  ;
        ANTENNAGATEAREA 0.372  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.020 5.500 1.220 ;
        LAYER ME2 ;
        RECT  5.300 0.800 5.500 1.350 ;
        LAYER ME1 ;
        RECT  5.120 1.020 6.120 1.220 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.540 1.470 10.740 2.540 ;
        RECT  9.500 1.840 9.700 2.540 ;
        RECT  8.460 1.840 8.660 2.540 ;
        RECT  7.420 1.840 7.620 2.540 ;
        RECT  6.380 1.480 6.580 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.540 -0.140 10.740 0.660 ;
        RECT  9.460 -0.140 9.740 0.500 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 1.480 2.980 1.680 ;
        RECT  1.700 1.480 1.900 2.080 ;
        RECT  3.260 1.520 4.540 1.720 ;
        RECT  3.260 1.520 3.460 2.080 ;
        RECT  2.180 1.880 3.460 2.080 ;
        RECT  4.820 1.440 6.060 1.640 ;
        RECT  4.820 1.440 5.020 2.080 ;
        RECT  3.740 1.880 5.020 2.080 ;
        RECT  5.860 1.440 6.060 2.080 ;
        RECT  0.660 0.380 0.860 0.820 ;
        RECT  1.700 0.380 1.900 0.820 ;
        RECT  2.740 0.380 2.940 0.820 ;
        RECT  3.780 0.380 3.980 0.820 ;
        RECT  4.820 0.380 5.020 0.820 ;
        RECT  5.860 0.380 6.060 0.820 ;
        RECT  0.140 0.660 6.580 0.820 ;
        RECT  6.380 0.660 6.580 1.220 ;
        RECT  6.380 1.020 8.040 1.220 ;
        RECT  0.140 0.660 0.340 2.080 ;
        RECT  0.140 1.880 1.420 2.080 ;
        RECT  9.080 1.020 10.440 1.220 ;
        LAYER VTPH ;
        RECT  0.000 1.140 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
    END
END OR4M16HM

MACRO OR4M12HM
    CLASS CORE ;
    FOREIGN OR4M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.379  LAYER ME1  ;
        ANTENNAGATEAREA 0.379  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.646  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.020 2.300 1.220 ;
        LAYER ME2 ;
        RECT  2.100 0.800 2.300 1.350 ;
        LAYER ME1 ;
        RECT  2.000 1.020 3.000 1.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.379  LAYER ME1  ;
        ANTENNAGATEAREA 0.379  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.646  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.800 1.100 1.350 ;
        LAYER ME1 ;
        RECT  0.500 1.020 1.500 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.416  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.980 0.380 9.180 2.080 ;
        RECT  6.900 1.440 9.180 1.640 ;
        RECT  8.850 0.660 9.180 1.640 ;
        RECT  6.900 0.660 9.180 0.860 ;
        RECT  7.940 1.440 8.140 2.080 ;
        RECT  7.940 0.380 8.140 0.860 ;
        RECT  6.900 1.440 7.100 2.080 ;
        RECT  6.900 0.380 7.100 0.860 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.379  LAYER ME1  ;
        ANTENNAGATEAREA 0.379  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.646  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.020 3.900 1.220 ;
        LAYER ME2 ;
        RECT  3.700 0.800 3.900 1.350 ;
        LAYER ME1 ;
        RECT  3.560 1.020 4.560 1.220 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.379  LAYER ME1  ;
        ANTENNAGATEAREA 0.379  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.646  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.020 5.500 1.220 ;
        LAYER ME2 ;
        RECT  5.300 0.800 5.500 1.350 ;
        LAYER ME1 ;
        RECT  5.120 1.020 6.120 1.220 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.500 1.480 9.700 2.540 ;
        RECT  8.460 1.840 8.660 2.540 ;
        RECT  7.420 1.840 7.620 2.540 ;
        RECT  6.380 1.480 6.580 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.500 -0.140 9.700 0.660 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 1.480 2.980 1.680 ;
        RECT  1.700 1.480 1.900 2.080 ;
        RECT  3.260 1.520 4.540 1.720 ;
        RECT  3.260 1.520 3.460 2.080 ;
        RECT  2.180 1.880 3.460 2.080 ;
        RECT  4.820 1.440 6.060 1.640 ;
        RECT  4.820 1.440 5.020 2.080 ;
        RECT  3.740 1.880 5.020 2.080 ;
        RECT  5.860 1.440 6.060 2.080 ;
        RECT  0.660 0.380 0.860 0.820 ;
        RECT  1.700 0.380 1.900 0.820 ;
        RECT  2.740 0.380 2.940 0.820 ;
        RECT  3.780 0.380 3.980 0.820 ;
        RECT  4.820 0.380 5.020 0.820 ;
        RECT  5.860 0.380 6.060 0.820 ;
        RECT  0.140 0.660 6.580 0.820 ;
        RECT  6.380 0.660 6.580 1.220 ;
        RECT  6.380 1.020 8.400 1.220 ;
        RECT  0.140 0.660 0.340 2.080 ;
        RECT  0.140 1.880 1.420 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
    END
END OR4M12HM

MACRO OR4M0HM
    CLASS CORE ;
    FOREIGN OR4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.100 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.080 1.100 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.080 1.680 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.880 1.080 2.300 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 0.340 3.100 1.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.100 2.080 2.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.300 -0.140 2.580 0.540 ;
        RECT  1.180 -0.140 1.460 0.540 ;
        RECT  0.140 -0.140 0.340 0.840 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.610 0.620 0.900 0.920 ;
        RECT  1.740 0.620 2.020 0.920 ;
        RECT  0.610 0.760 2.640 0.920 ;
        RECT  2.460 0.760 2.640 1.920 ;
        RECT  0.100 1.720 2.640 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OR4M0HM

MACRO OR3M8HM
    CLASS CORE ;
    FOREIGN OR3M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.520  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.160 1.050 2.360 1.250 ;
        LAYER ME2 ;
        RECT  2.100 0.950 2.360 1.560 ;
        LAYER ME1 ;
        RECT  2.160 0.980 2.420 1.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.620 2.840 1.780 ;
        RECT  2.640 0.990 2.840 1.780 ;
        RECT  1.300 0.990 1.500 1.780 ;
        RECT  1.000 0.990 1.500 1.270 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.070 1.030 3.400 1.230 ;
        RECT  0.500 1.940 3.270 2.100 ;
        RECT  3.070 1.030 3.270 2.100 ;
        RECT  0.500 0.990 0.700 2.100 ;
        RECT  0.320 0.990 0.700 1.270 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.130 1.440 5.330 2.080 ;
        RECT  4.090 0.680 5.330 0.860 ;
        RECT  5.130 0.430 5.330 0.860 ;
        RECT  4.090 1.440 5.330 1.640 ;
        RECT  4.900 0.680 5.100 1.640 ;
        RECT  4.090 1.440 4.290 2.080 ;
        RECT  4.090 0.430 4.290 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.650 1.450 5.850 2.540 ;
        RECT  4.570 1.870 4.850 2.540 ;
        RECT  3.500 1.450 3.780 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.650 -0.140 5.850 0.710 ;
        RECT  4.570 -0.140 4.850 0.500 ;
        RECT  3.460 -0.140 3.740 0.500 ;
        RECT  2.260 -0.140 2.540 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.340 0.860 0.820 ;
        RECT  1.700 0.340 1.900 1.460 ;
        RECT  2.820 0.310 3.020 0.820 ;
        RECT  0.660 0.660 3.720 0.820 ;
        RECT  3.560 0.660 3.720 1.240 ;
        RECT  3.560 1.040 4.510 1.240 ;
        RECT  1.700 0.660 1.980 1.460 ;
        LAYER VTPH ;
        RECT  1.320 0.940 2.420 2.400 ;
        RECT  0.000 1.100 3.520 2.400 ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 0.940 ;
        RECT  0.000 0.000 1.320 1.100 ;
        RECT  2.420 0.000 6.000 1.100 ;
        RECT  3.520 0.000 6.000 1.140 ;
    END
END OR3M8HM

MACRO OR3M6HM
    CLASS CORE ;
    FOREIGN OR3M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        ANTENNAGATEAREA 0.212  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.154  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.340 1.180 1.540 1.380 ;
        LAYER ME2 ;
        RECT  1.300 1.120 1.560 1.560 ;
        LAYER ME1 ;
        RECT  1.280 1.120 1.880 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.580 2.320 1.740 ;
        RECT  2.120 1.150 2.320 1.740 ;
        RECT  0.800 1.120 1.100 1.740 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.800 2.900 1.340 ;
        RECT  0.320 0.800 2.900 0.960 ;
        RECT  0.320 0.800 0.520 1.320 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.460 0.430 4.700 2.080 ;
        RECT  3.420 1.440 4.700 1.640 ;
        RECT  3.420 0.680 4.700 0.860 ;
        RECT  3.420 1.440 3.620 2.080 ;
        RECT  3.420 0.430 3.620 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.900 1.870 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        RECT  0.140 1.680 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.900 -0.140 4.180 0.500 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        RECT  1.700 -0.140 1.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.100 0.480 3.220 0.640 ;
        RECT  3.060 0.480 3.220 1.700 ;
        RECT  3.060 1.040 4.270 1.240 ;
        RECT  3.060 1.040 3.230 1.700 ;
        RECT  2.480 1.540 3.230 1.700 ;
        RECT  2.480 1.540 2.640 2.060 ;
        RECT  1.380 1.900 2.640 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OR3M6HM

MACRO OR3M4HM
    CLASS CORE ;
    FOREIGN OR3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.020 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.020 1.700 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 1.440 2.700 1.640 ;
        RECT  2.500 0.720 2.700 1.640 ;
        RECT  2.220 0.720 2.700 0.920 ;
        RECT  2.220 1.440 2.420 2.080 ;
        RECT  2.220 0.390 2.420 0.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.740 1.840 2.940 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.740 -0.140 2.940 0.560 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.340 1.380 0.820 ;
        RECT  0.140 0.660 2.020 0.820 ;
        RECT  1.860 0.660 2.020 1.280 ;
        RECT  1.860 1.080 2.280 1.280 ;
        RECT  0.140 0.340 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OR3M4HM

MACRO OR3M2HM
    CLASS CORE ;
    FOREIGN OR3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.020 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.300 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.020 1.900 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.292  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.330 2.700 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.930 1.840 2.130 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.400 1.540 0.820 ;
        RECT  0.140 0.660 2.300 0.820 ;
        RECT  2.140 0.660 2.300 1.360 ;
        RECT  0.140 0.420 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OR3M2HM

MACRO OR3M1HM
    CLASS CORE ;
    FOREIGN OR3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.020 0.700 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.300 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.020 1.900 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.320 2.700 2.000 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.930 1.840 2.130 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.400 1.540 0.820 ;
        RECT  0.140 0.660 2.300 0.820 ;
        RECT  2.140 0.660 2.300 1.360 ;
        RECT  0.140 0.420 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OR3M1HM

MACRO OR3M16HM
    CLASS CORE ;
    FOREIGN OR3M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.020 2.700 1.220 ;
        LAYER ME2 ;
        RECT  2.500 0.800 2.700 1.350 ;
        LAYER ME1 ;
        RECT  2.260 1.020 3.260 1.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.181  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.800 1.100 1.350 ;
        LAYER ME1 ;
        RECT  0.700 1.020 1.350 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.888  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.720 1.440 8.920 2.080 ;
        RECT  5.600 0.660 8.920 0.860 ;
        RECT  8.720 0.380 8.920 0.860 ;
        RECT  5.600 1.440 8.920 1.630 ;
        RECT  7.680 1.440 7.880 2.080 ;
        RECT  7.680 0.380 7.880 0.860 ;
        RECT  5.600 1.440 7.880 1.640 ;
        RECT  7.250 0.660 7.550 1.640 ;
        RECT  6.640 1.440 6.840 2.080 ;
        RECT  6.640 0.380 6.840 0.860 ;
        RECT  5.600 1.440 5.800 2.080 ;
        RECT  5.600 0.380 5.800 0.860 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        ANTENNAGATEAREA 0.374  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.020 4.300 1.220 ;
        LAYER ME2 ;
        RECT  4.100 0.800 4.300 1.350 ;
        LAYER ME1 ;
        RECT  3.820 1.020 4.820 1.220 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.240 1.470 9.440 2.540 ;
        RECT  8.200 1.840 8.400 2.540 ;
        RECT  7.160 1.840 7.360 2.540 ;
        RECT  6.120 1.840 6.320 2.540 ;
        RECT  5.080 1.480 5.280 2.540 ;
        RECT  4.040 1.840 4.240 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.240 -0.140 9.440 0.660 ;
        RECT  8.160 -0.140 8.440 0.500 ;
        RECT  7.120 -0.140 7.400 0.500 ;
        RECT  6.080 -0.140 6.360 0.500 ;
        RECT  5.040 -0.140 5.320 0.500 ;
        RECT  4.000 -0.140 4.280 0.500 ;
        RECT  2.960 -0.140 3.240 0.500 ;
        RECT  1.920 -0.140 2.200 0.500 ;
        RECT  0.880 -0.140 1.160 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.960 1.520 3.240 1.720 ;
        RECT  1.960 1.520 2.160 2.080 ;
        RECT  0.880 1.880 2.160 2.080 ;
        RECT  3.520 1.440 4.760 1.640 ;
        RECT  3.520 1.440 3.720 2.080 ;
        RECT  2.440 1.880 3.720 2.080 ;
        RECT  4.560 1.440 4.760 2.080 ;
        RECT  0.400 0.380 0.600 0.820 ;
        RECT  1.440 0.380 1.640 0.820 ;
        RECT  2.480 0.380 2.680 0.820 ;
        RECT  3.520 0.380 3.720 0.820 ;
        RECT  4.560 0.380 4.760 0.820 ;
        RECT  0.400 0.660 5.280 0.820 ;
        RECT  5.080 0.660 5.280 1.220 ;
        RECT  5.080 1.020 6.740 1.220 ;
        RECT  1.510 0.660 1.710 1.680 ;
        RECT  0.400 1.480 1.710 1.680 ;
        RECT  0.400 1.480 0.600 2.080 ;
        RECT  7.780 1.020 9.140 1.220 ;
        LAYER VTPH ;
        RECT  0.000 1.080 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.080 ;
    END
END OR3M16HM

MACRO OR3M12HM
    CLASS CORE ;
    FOREIGN OR3M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.364  LAYER ME1  ;
        ANTENNAGATEAREA 0.364  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.216  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.640 1.020 0.840 1.220 ;
        LAYER ME2 ;
        RECT  0.500 0.800 0.840 1.350 ;
        LAYER ME1 ;
        RECT  0.440 1.020 1.090 1.220 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.364  LAYER ME1  ;
        ANTENNAGATEAREA 0.364  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.716  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.020 2.300 1.220 ;
        LAYER ME2 ;
        RECT  2.100 0.800 2.300 1.350 ;
        LAYER ME1 ;
        RECT  2.000 1.020 3.000 1.220 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.420 1.440 7.620 2.080 ;
        RECT  5.340 0.660 7.620 0.860 ;
        RECT  7.420 0.380 7.620 0.860 ;
        RECT  5.340 1.440 7.620 1.640 ;
        RECT  6.440 0.660 6.740 1.640 ;
        RECT  6.380 1.440 6.580 2.080 ;
        RECT  6.380 0.380 6.580 0.860 ;
        RECT  5.340 1.440 5.540 2.080 ;
        RECT  5.340 0.380 5.540 0.860 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.364  LAYER ME1  ;
        ANTENNAGATEAREA 0.364  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.716  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.020 3.900 1.220 ;
        LAYER ME2 ;
        RECT  3.700 0.800 3.900 1.350 ;
        LAYER ME1 ;
        RECT  3.560 1.020 4.560 1.220 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.940 1.450 8.140 2.540 ;
        RECT  6.900 1.840 7.100 2.540 ;
        RECT  5.860 1.840 6.060 2.540 ;
        RECT  4.820 1.800 5.020 2.540 ;
        RECT  3.780 1.840 3.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.900 -0.140 8.180 0.500 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.700 1.520 2.980 1.720 ;
        RECT  1.700 1.520 1.900 2.080 ;
        RECT  0.620 1.880 1.900 2.080 ;
        RECT  3.260 1.440 4.500 1.640 ;
        RECT  3.260 1.440 3.460 2.080 ;
        RECT  2.180 1.880 3.460 2.080 ;
        RECT  4.300 1.440 4.500 2.080 ;
        RECT  0.140 0.300 0.340 0.820 ;
        RECT  1.180 0.300 1.380 0.820 ;
        RECT  2.220 0.300 2.420 0.820 ;
        RECT  3.260 0.300 3.460 0.820 ;
        RECT  4.300 0.300 4.500 0.820 ;
        RECT  0.140 0.660 5.020 0.820 ;
        RECT  4.820 0.660 5.020 1.220 ;
        RECT  4.820 1.020 6.180 1.220 ;
        RECT  1.250 0.660 1.450 1.680 ;
        RECT  0.140 1.480 1.450 1.680 ;
        RECT  0.140 1.480 0.340 2.080 ;
        RECT  6.920 1.020 7.780 1.220 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END OR3M12HM

MACRO OR3M0HM
    CLASS CORE ;
    FOREIGN OR3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.080 0.720 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.180 1.300 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.080 1.900 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.310 2.700 2.020 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.930 1.840 2.130 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.310 1.540 0.820 ;
        RECT  0.140 0.660 2.300 0.820 ;
        RECT  2.140 0.660 2.300 1.360 ;
        RECT  0.140 0.310 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OR3M0HM

MACRO OR2M8HM
    CLASS CORE ;
    FOREIGN OR2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        ANTENNAGATEAREA 0.252  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.816  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.810 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 1.020 1.600 1.260 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 2.060 1.600 ;
        RECT  1.860 1.000 2.060 1.600 ;
        RECT  0.500 1.000 0.700 1.600 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.976  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.800 0.410 4.020 2.090 ;
        RECT  2.740 1.500 4.020 1.660 ;
        RECT  3.700 0.680 4.020 1.660 ;
        RECT  2.740 0.680 4.020 0.880 ;
        RECT  2.740 1.500 2.940 2.020 ;
        RECT  2.740 0.410 2.940 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.300 1.480 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.080 2.080 2.360 2.540 ;
        RECT  0.340 1.840 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.300 -0.140 4.500 0.690 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.340 0.860 0.840 ;
        RECT  1.700 0.340 1.900 0.840 ;
        RECT  0.660 0.680 2.460 0.840 ;
        RECT  2.300 1.080 3.540 1.280 ;
        RECT  2.300 0.680 2.460 1.920 ;
        RECT  1.100 1.760 2.460 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OR2M8HM

MACRO OR2M6HM
    CLASS CORE ;
    FOREIGN OR2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.560 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.820 1.000 1.100 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.903  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 1.540 3.100 2.090 ;
        RECT  2.900 0.410 3.100 2.090 ;
        RECT  1.700 0.680 3.100 0.880 ;
        RECT  2.760 0.410 3.100 0.880 ;
        RECT  1.660 1.540 3.100 1.740 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  1.660 1.540 1.880 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.040 2.080 1.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.100 -0.140 0.380 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.300 0.840 0.840 ;
        RECT  0.680 0.680 1.420 0.840 ;
        RECT  1.260 1.080 2.500 1.280 ;
        RECT  1.260 0.680 1.420 1.920 ;
        RECT  0.100 1.720 1.420 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OR2M6HM

MACRO OR2M4HM
    CLASS CORE ;
    FOREIGN OR2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.500 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.000 1.100 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.540 2.700 1.740 ;
        RECT  2.490 0.680 2.700 1.740 ;
        RECT  1.640 0.680 2.700 0.880 ;
        RECT  1.640 0.360 1.960 0.880 ;
        RECT  1.640 1.540 1.950 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.040 2.080 1.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.100 -0.140 0.380 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.300 0.840 0.840 ;
        RECT  0.680 0.680 1.420 0.840 ;
        RECT  1.260 1.080 2.120 1.280 ;
        RECT  1.260 0.680 1.420 1.920 ;
        RECT  0.100 1.720 1.420 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OR2M4HM

MACRO OR2M2HM
    CLASS CORE ;
    FOREIGN OR2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 0.600 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.040 1.140 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.450 1.900 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.040 2.080 1.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.100 -0.140 1.300 0.380 ;
        RECT  0.140 -0.140 0.340 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.560 1.500 0.880 ;
        RECT  1.300 0.560 1.500 1.920 ;
        RECT  0.180 1.760 1.500 1.920 ;
        RECT  0.180 1.760 0.380 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END OR2M2HM

MACRO OR2M1HM
    CLASS CORE ;
    FOREIGN OR2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 0.600 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.040 1.140 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.450 1.900 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.040 2.080 1.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.100 -0.140 1.300 0.380 ;
        RECT  0.140 -0.140 0.340 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.560 1.500 0.880 ;
        RECT  1.300 0.560 1.500 1.920 ;
        RECT  0.180 1.760 1.500 1.920 ;
        RECT  0.180 1.760 0.380 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END OR2M1HM

MACRO OR2M16HM
    CLASS CORE ;
    FOREIGN OR2M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.370  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.800 0.800 2.420 1.270 ;
        RECT  0.460 0.800 2.420 0.960 ;
        RECT  0.460 0.800 0.710 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.370  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.440 2.860 1.600 ;
        RECT  2.620 1.000 2.860 1.600 ;
        RECT  0.900 1.120 1.280 1.600 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.600 1.510 6.820 2.100 ;
        RECT  3.460 0.680 6.780 0.840 ;
        RECT  6.580 0.370 6.780 0.840 ;
        RECT  3.420 1.510 6.820 1.710 ;
        RECT  5.540 0.660 6.780 0.840 ;
        RECT  5.540 1.510 5.740 2.100 ;
        RECT  5.540 0.370 5.740 0.840 ;
        RECT  4.900 0.680 5.500 1.710 ;
        RECT  4.500 1.510 4.700 2.100 ;
        RECT  4.500 0.370 4.700 0.840 ;
        RECT  3.460 0.370 3.660 0.840 ;
        RECT  3.420 1.510 3.640 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  7.060 1.900 7.340 2.540 ;
        RECT  6.020 1.900 6.300 2.540 ;
        RECT  4.980 1.900 5.260 2.540 ;
        RECT  3.940 1.900 4.220 2.540 ;
        RECT  2.860 2.080 3.140 2.540 ;
        RECT  1.100 2.080 1.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.060 -0.140 7.340 0.500 ;
        RECT  6.020 -0.140 6.300 0.500 ;
        RECT  4.980 -0.140 5.260 0.500 ;
        RECT  3.940 -0.140 4.220 0.520 ;
        RECT  2.860 -0.140 3.140 0.320 ;
        RECT  1.740 -0.140 2.020 0.320 ;
        RECT  0.700 -0.140 0.900 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.480 3.200 0.640 ;
        RECT  3.040 1.040 4.740 1.240 ;
        RECT  3.040 0.480 3.200 1.920 ;
        RECT  0.180 1.760 3.200 1.920 ;
        RECT  5.660 1.040 7.010 1.240 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END OR2M16HM

MACRO OR2M12HM
    CLASS CORE ;
    FOREIGN OR2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.370  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.800 0.800 2.420 1.270 ;
        RECT  0.460 0.800 2.420 0.960 ;
        RECT  0.460 0.800 0.710 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.440 2.860 1.600 ;
        RECT  2.620 1.000 2.860 1.600 ;
        RECT  0.900 1.120 1.280 1.600 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.540 1.510 5.780 2.100 ;
        RECT  3.460 0.680 5.740 0.840 ;
        RECT  5.540 0.370 5.740 0.840 ;
        RECT  3.420 1.510 5.780 1.710 ;
        RECT  4.900 0.680 5.500 1.710 ;
        RECT  4.500 1.510 4.700 2.100 ;
        RECT  4.500 0.370 4.700 0.840 ;
        RECT  3.460 0.370 3.660 0.840 ;
        RECT  3.420 1.510 3.640 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  6.020 1.900 6.300 2.540 ;
        RECT  4.980 1.900 5.260 2.540 ;
        RECT  3.940 1.900 4.220 2.540 ;
        RECT  2.860 2.080 3.140 2.540 ;
        RECT  1.100 2.080 1.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  6.020 -0.140 6.300 0.500 ;
        RECT  4.980 -0.140 5.260 0.500 ;
        RECT  3.940 -0.140 4.220 0.520 ;
        RECT  2.860 -0.140 3.140 0.320 ;
        RECT  1.740 -0.140 2.020 0.320 ;
        RECT  0.700 -0.140 0.900 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.480 3.200 0.640 ;
        RECT  3.040 1.040 4.740 1.240 ;
        RECT  3.040 0.480 3.200 1.920 ;
        RECT  0.180 1.760 3.200 1.920 ;
        RECT  5.660 1.040 6.240 1.240 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END OR2M12HM

MACRO OR2M0HM
    CLASS CORE ;
    FOREIGN OR2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 0.600 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.040 1.140 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.450 1.900 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.040 2.080 1.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.100 -0.140 1.300 0.380 ;
        RECT  0.140 -0.140 0.340 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.560 1.500 0.880 ;
        RECT  1.300 0.560 1.500 1.920 ;
        RECT  0.180 1.760 1.500 1.920 ;
        RECT  0.180 1.760 0.380 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END OR2M0HM

MACRO OAI33M8HM
    CLASS CORE ;
    FOREIGN OAI33M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.523  LAYER ME1  ;
        ANTENNAGATEAREA 0.523  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.729  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.100 1.040 10.300 1.240 ;
        LAYER ME2 ;
        RECT  10.100 0.840 10.300 1.560 ;
        LAYER ME1 ;
        RECT  9.820 1.040 11.340 1.260 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        ANTENNAGATEAREA 0.504  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.754  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.040 8.300 1.240 ;
        LAYER ME2 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  7.260 1.040 8.740 1.260 ;
        END
    END A1
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.514  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 2.100 1.240 ;
        RECT  0.100 0.840 0.300 1.240 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.625  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.450 0.620 13.230 0.780 ;
        RECT  4.820 1.580 9.260 1.740 ;
        RECT  8.900 1.540 9.260 1.740 ;
        RECT  8.900 0.620 9.100 1.740 ;
        RECT  4.820 1.540 5.110 1.740 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        ANTENNAGATEAREA 0.528  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.842  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  12.100 1.040 12.300 1.240 ;
        LAYER ME2 ;
        RECT  12.100 0.840 12.300 1.560 ;
        LAYER ME1 ;
        RECT  11.880 1.040 13.530 1.260 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.514  LAYER ME1  ;
        ANTENNAGATEAREA 0.514  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.701  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.040 6.300 1.240 ;
        LAYER ME2 ;
        RECT  6.100 0.840 6.300 1.560 ;
        LAYER ME1 ;
        RECT  5.260 1.040 6.740 1.240 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.514  LAYER ME1  ;
        ANTENNAGATEAREA 0.514  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.701  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.700 1.040 4.180 1.240 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.100 1.900 13.380 2.540 ;
        RECT  12.060 1.900 12.340 2.540 ;
        RECT  1.740 1.900 2.020 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  6.320 -0.140 6.630 0.460 ;
        RECT  5.210 -0.140 5.500 0.460 ;
        RECT  3.960 -0.140 4.240 0.460 ;
        RECT  2.820 -0.140 3.100 0.460 ;
        RECT  1.650 -0.140 1.930 0.460 ;
        RECT  0.450 -0.140 0.730 0.460 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 1.480 4.620 1.640 ;
        RECT  2.300 1.480 4.620 1.680 ;
        RECT  0.180 1.480 0.400 2.100 ;
        RECT  1.260 1.480 1.460 2.100 ;
        RECT  2.300 1.480 2.500 2.100 ;
        RECT  2.750 1.860 4.160 2.060 ;
        RECT  2.750 1.900 6.710 2.060 ;
        RECT  7.350 1.900 11.370 2.060 ;
        RECT  6.940 0.300 13.650 0.460 ;
        RECT  1.080 0.380 1.280 0.800 ;
        RECT  2.300 0.380 2.500 0.800 ;
        RECT  3.440 0.380 3.640 0.800 ;
        RECT  5.810 0.380 6.010 0.800 ;
        RECT  13.490 0.300 13.650 0.760 ;
        RECT  6.940 0.300 7.140 0.800 ;
        RECT  1.080 0.640 7.140 0.800 ;
        RECT  9.420 1.580 13.900 1.740 ;
        RECT  13.600 1.580 13.900 1.780 ;
        LAYER VTPH ;
        RECT  9.280 1.100 10.160 2.400 ;
        RECT  0.000 1.140 7.340 2.400 ;
        RECT  9.280 1.140 14.000 2.400 ;
        RECT  0.000 1.160 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.100 ;
        RECT  0.000 0.000 9.280 1.140 ;
        RECT  10.160 0.000 14.000 1.140 ;
        RECT  7.340 0.000 9.280 1.160 ;
    END
END OAI33M8HM

MACRO OAI33M4HM
    CLASS CORE ;
    FOREIGN OAI33M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.257  LAYER ME1  ;
        ANTENNAGATEAREA 0.257  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.924  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.070 2.700 1.270 ;
        LAYER ME2 ;
        RECT  2.500 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.320 1.030 2.920 1.380 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        ANTENNAGATEAREA 0.278  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.718  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.080 5.500 1.280 ;
        LAYER ME2 ;
        RECT  5.300 0.980 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.200 1.080 5.920 1.280 ;
        END
    END A3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        ANTENNAGATEAREA 0.278  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.513  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.350 1.080 3.550 1.280 ;
        LAYER ME2 ;
        RECT  3.300 0.950 3.550 1.560 ;
        LAYER ME1 ;
        RECT  3.250 1.080 3.860 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.720 1.440 6.360 1.600 ;
        RECT  6.100 1.060 6.360 1.600 ;
        RECT  4.720 1.060 4.920 1.600 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.257  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.440 2.040 1.600 ;
        RECT  1.840 1.020 2.040 1.600 ;
        RECT  0.280 1.100 0.700 1.600 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.740 0.740 6.180 0.900 ;
        RECT  5.900 0.620 6.180 0.900 ;
        RECT  4.860 0.620 5.140 0.900 ;
        RECT  2.460 1.540 4.340 1.700 ;
        RECT  4.100 0.740 4.340 1.700 ;
        RECT  3.740 0.620 4.020 0.900 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.257  LAYER ME1  ;
        ANTENNAGATEAREA 0.257  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.863  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.830 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 1.000 1.600 1.280 ;
        END
    END B3
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.420 2.080 5.700 2.540 ;
        RECT  1.040 2.080 1.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.760 2.220 1.920 ;
        RECT  0.140 1.760 0.340 2.040 ;
        RECT  2.020 1.900 3.340 2.060 ;
        RECT  4.580 1.760 6.620 1.920 ;
        RECT  3.500 1.860 4.780 2.060 ;
        RECT  3.280 0.300 6.660 0.460 ;
        RECT  4.300 0.300 4.580 0.580 ;
        RECT  5.380 0.300 5.660 0.580 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  2.220 0.380 2.420 0.820 ;
        RECT  6.460 0.300 6.660 0.760 ;
        RECT  3.280 0.300 3.440 0.820 ;
        RECT  0.140 0.660 3.440 0.820 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END OAI33M4HM

MACRO OAI33M2HM
    CLASS CORE ;
    FOREIGN OAI33M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.100 1.120 1.560 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.500 1.560 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.095  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.030 1.220 2.230 1.420 ;
        LAYER ME2 ;
        RECT  2.030 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.940 1.100 2.280 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.100 2.720 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 1.100 3.200 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.100 1.600 1.560 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.774  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.690 1.740 3.520 1.900 ;
        RECT  3.360 0.300 3.520 1.900 ;
        RECT  3.200 0.300 3.520 0.840 ;
        RECT  2.180 0.300 3.520 0.460 ;
        RECT  2.180 0.300 2.460 0.620 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 2.080 3.500 2.540 ;
        RECT  0.180 1.840 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  1.140 -0.140 1.420 0.620 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.420 0.840 0.940 ;
        RECT  1.720 0.410 1.880 0.940 ;
        RECT  2.700 0.620 2.980 0.940 ;
        RECT  0.680 0.780 2.980 0.940 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI33M2HM

MACRO OAI33M1HM
    CLASS CORE ;
    FOREIGN OAI33M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.100 1.120 1.560 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.500 1.560 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        ANTENNAGATEAREA 0.096  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.000 1.180 2.200 1.380 ;
        LAYER ME2 ;
        RECT  2.000 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.940 1.100 2.280 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.100 2.720 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 1.100 3.200 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.100 1.600 1.560 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.874  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.690 1.740 3.520 1.900 ;
        RECT  3.360 0.300 3.520 1.900 ;
        RECT  3.200 0.300 3.520 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 2.080 3.500 2.540 ;
        RECT  0.180 1.840 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  1.140 -0.140 1.420 0.620 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.390 0.840 0.940 ;
        RECT  1.720 0.390 1.880 0.940 ;
        RECT  2.760 0.520 2.920 0.940 ;
        RECT  0.680 0.780 2.920 0.940 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI33M1HM

MACRO OAI33M0HM
    CLASS CORE ;
    FOREIGN OAI33M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.100 1.120 1.560 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.500 1.560 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.253  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.030 1.230 2.230 1.430 ;
        LAYER ME2 ;
        RECT  2.030 0.830 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.940 1.100 2.280 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.100 2.720 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 1.100 3.200 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.100 1.600 1.560 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.795  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.690 1.740 3.520 1.900 ;
        RECT  3.360 0.300 3.520 1.900 ;
        RECT  3.200 0.300 3.520 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 2.080 3.500 2.540 ;
        RECT  0.180 1.790 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  1.140 -0.140 1.420 0.620 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.360 0.840 0.940 ;
        RECT  1.720 0.360 1.880 0.940 ;
        RECT  2.760 0.520 2.920 0.940 ;
        RECT  0.680 0.780 2.920 0.940 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI33M0HM

MACRO OAI32M8HM
    CLASS CORE ;
    FOREIGN OAI32M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        ANTENNAGATEAREA 0.528  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.655  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.020 3.500 1.220 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.620 1.020 4.100 1.220 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        ANTENNAGATEAREA 0.528  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.389  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.020 6.300 1.220 ;
        LAYER ME2 ;
        RECT  6.100 0.840 6.300 1.560 ;
        LAYER ME1 ;
        RECT  5.490 1.020 6.700 1.220 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 2.060 1.180 ;
        RECT  0.100 0.840 0.840 1.180 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.860 1.930 8.140 2.100 ;
        RECT  7.860 1.900 8.140 2.100 ;
        RECT  6.860 1.500 7.060 2.100 ;
        RECT  4.700 1.500 7.060 1.660 ;
        RECT  1.140 0.700 6.580 0.860 ;
        RECT  6.300 0.620 6.580 0.860 ;
        RECT  4.860 0.620 5.540 0.860 ;
        RECT  4.900 0.620 5.100 1.660 ;
        RECT  3.220 0.620 3.500 0.860 ;
        RECT  2.180 0.620 2.460 0.860 ;
        RECT  1.140 0.620 1.420 0.860 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.004  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.700 1.020 7.900 1.220 ;
        LAYER ME2 ;
        RECT  7.700 0.840 7.900 1.560 ;
        LAYER ME1 ;
        RECT  7.160 1.020 8.660 1.240 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.561  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.700 1.020 9.900 1.220 ;
        LAYER ME2 ;
        RECT  9.700 0.840 9.900 1.560 ;
        LAYER ME1 ;
        RECT  9.240 1.020 10.360 1.240 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  9.900 1.900 10.180 2.540 ;
        RECT  8.860 1.900 9.140 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  9.900 -0.140 10.180 0.540 ;
        RECT  8.860 -0.140 9.140 0.540 ;
        RECT  7.340 -0.140 7.620 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.460 4.540 1.660 ;
        RECT  0.100 1.460 0.320 2.080 ;
        RECT  1.180 1.460 1.380 2.080 ;
        RECT  2.220 1.460 2.420 2.080 ;
        RECT  2.660 1.900 6.620 2.060 ;
        RECT  7.340 1.500 10.660 1.660 ;
        RECT  7.340 1.500 7.620 1.770 ;
        RECT  8.380 1.500 8.660 1.770 ;
        RECT  9.420 1.500 9.620 2.000 ;
        RECT  10.460 1.500 10.660 2.000 ;
        RECT  0.620 0.300 7.060 0.460 ;
        RECT  0.620 0.300 0.900 0.540 ;
        RECT  1.660 0.300 1.940 0.540 ;
        RECT  2.700 0.300 2.980 0.540 ;
        RECT  3.740 0.300 4.020 0.540 ;
        RECT  5.780 0.300 6.060 0.540 ;
        RECT  6.860 0.300 7.060 0.860 ;
        RECT  7.900 0.480 8.100 0.860 ;
        RECT  9.380 0.480 9.660 0.860 ;
        RECT  10.460 0.480 10.660 0.860 ;
        RECT  6.860 0.700 10.660 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.800 1.140 ;
    END
END OAI32M8HM

MACRO OAI32M4HM
    CLASS CORE ;
    FOREIGN OAI32M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME2  ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.420  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.060 2.700 1.260 ;
        LAYER ME1 ;
        RECT  2.440 1.060 3.000 1.260 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.360 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.960 1.440 5.540 1.600 ;
        RECT  5.300 1.060 5.540 1.600 ;
        RECT  3.960 1.060 4.160 1.600 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 2.280 1.600 ;
        RECT  2.080 1.060 2.280 1.600 ;
        RECT  0.500 1.060 0.860 1.600 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.256  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.940 0.740 5.380 0.900 ;
        RECT  5.100 0.620 5.380 0.900 ;
        RECT  4.060 0.620 4.340 0.900 ;
        RECT  3.300 0.740 3.500 1.780 ;
        RECT  2.460 1.440 3.500 1.600 ;
        RECT  2.940 0.620 3.220 0.900 ;
        RECT  0.420 1.760 2.620 1.920 ;
        RECT  2.460 1.440 2.620 1.920 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        ANTENNAGATEAREA 0.278  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.569  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.060 4.700 1.260 ;
        LAYER ME1 ;
        RECT  4.440 1.060 5.080 1.260 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.360 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        ANTENNAGATEAREA 0.252  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.733  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.060 1.500 1.260 ;
        LAYER ME1 ;
        RECT  1.200 1.060 1.840 1.260 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.360 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  4.620 2.080 4.900 2.540 ;
        RECT  1.340 2.080 1.620 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  1.900 -0.140 2.180 0.580 ;
        RECT  0.860 -0.140 1.140 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.800 1.760 5.820 1.920 ;
        RECT  2.800 1.760 3.000 2.100 ;
        RECT  3.800 1.760 3.960 2.100 ;
        RECT  2.800 1.940 3.960 2.100 ;
        RECT  2.480 0.300 5.860 0.460 ;
        RECT  3.500 0.300 3.780 0.580 ;
        RECT  4.580 0.300 4.860 0.580 ;
        RECT  5.660 0.300 5.860 0.680 ;
        RECT  0.400 0.420 0.560 0.900 ;
        RECT  1.440 0.420 1.600 0.900 ;
        RECT  2.480 0.300 2.640 0.900 ;
        RECT  0.400 0.740 2.640 0.900 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END OAI32M4HM

MACRO OAI32M2HM
    CLASS CORE ;
    FOREIGN OAI32M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.020 1.650 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.330 1.700 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.010 1.020 2.370 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.020 3.100 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.646  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.540 1.780 2.090 1.940 ;
        RECT  0.100 0.700 1.470 0.860 ;
        RECT  1.190 0.620 1.470 0.860 ;
        RECT  0.540 0.700 0.740 1.940 ;
        RECT  0.100 0.440 0.380 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.750 1.900 3.030 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.230 -0.140 2.510 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.670 0.300 1.950 0.460 ;
        RECT  0.670 0.300 0.950 0.540 ;
        RECT  1.750 0.300 1.950 0.860 ;
        RECT  2.750 0.480 3.030 0.860 ;
        RECT  1.750 0.700 3.030 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI32M2HM

MACRO OAI32M1HM
    CLASS CORE ;
    FOREIGN OAI32M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.020 1.690 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.330 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.050 1.020 2.410 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.700 1.020 3.100 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.780 2.090 1.940 ;
        RECT  0.100 0.700 1.460 0.860 ;
        RECT  1.180 0.620 1.460 0.860 ;
        RECT  0.500 0.700 0.700 1.940 ;
        RECT  0.100 0.380 0.380 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.790 1.900 3.070 2.540 ;
        RECT  0.100 1.840 0.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.270 -0.140 2.550 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.300 1.990 0.460 ;
        RECT  0.620 0.300 0.900 0.540 ;
        RECT  1.790 0.300 1.990 0.860 ;
        RECT  2.790 0.320 3.070 0.860 ;
        RECT  1.790 0.700 3.070 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI32M1HM

MACRO OAI32M0HM
    CLASS CORE ;
    FOREIGN OAI32M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.020 1.690 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.330 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.050 1.020 2.410 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.700 1.020 3.100 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.900 2.130 2.060 ;
        RECT  0.100 0.700 1.460 0.860 ;
        RECT  1.180 0.620 1.460 0.860 ;
        RECT  0.500 0.700 0.700 2.060 ;
        RECT  0.100 0.380 0.380 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.790 1.900 3.070 2.540 ;
        RECT  0.100 1.840 0.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.270 -0.140 2.550 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.300 1.990 0.460 ;
        RECT  0.620 0.300 0.900 0.540 ;
        RECT  1.790 0.300 1.990 0.860 ;
        RECT  2.790 0.320 3.070 0.860 ;
        RECT  1.790 0.700 3.070 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI32M0HM

MACRO OAI31M8HM
    CLASS CORE ;
    FOREIGN OAI31M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        ANTENNAGATEAREA 0.528  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.655  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.020 3.500 1.220 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.660 1.020 4.140 1.220 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME2  ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.389  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.020 6.300 1.220 ;
        LAYER ME2 ;
        RECT  6.100 0.840 6.300 1.560 ;
        LAYER ME1 ;
        RECT  5.530 1.020 6.740 1.220 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.528  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 2.100 1.180 ;
        RECT  0.100 0.840 0.760 1.180 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.440 1.020 8.700 1.640 ;
        RECT  7.200 1.020 8.700 1.240 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.030  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.940 1.500 8.140 2.000 ;
        RECT  6.900 1.500 8.140 1.740 ;
        RECT  6.900 1.500 7.100 2.000 ;
        RECT  4.740 1.500 8.140 1.660 ;
        RECT  1.180 0.700 6.620 0.860 ;
        RECT  6.340 0.620 6.620 0.860 ;
        RECT  4.900 0.620 5.580 0.860 ;
        RECT  4.900 0.620 5.100 1.660 ;
        RECT  3.260 0.620 3.540 0.860 ;
        RECT  2.220 0.620 2.500 0.860 ;
        RECT  1.180 0.620 1.460 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  1.700 1.900 1.980 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.460 -0.140 8.660 0.760 ;
        RECT  7.380 -0.140 7.660 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.460 4.580 1.660 ;
        RECT  0.140 1.460 0.360 2.080 ;
        RECT  1.220 1.460 1.420 2.080 ;
        RECT  2.260 1.460 2.460 2.080 ;
        RECT  2.700 1.900 6.660 2.060 ;
        RECT  0.660 0.300 7.100 0.460 ;
        RECT  0.660 0.300 0.940 0.540 ;
        RECT  1.700 0.300 1.980 0.540 ;
        RECT  2.740 0.300 3.020 0.540 ;
        RECT  3.780 0.300 4.060 0.540 ;
        RECT  5.820 0.300 6.100 0.540 ;
        RECT  6.900 0.300 7.100 0.860 ;
        RECT  7.940 0.480 8.140 0.860 ;
        RECT  6.900 0.700 8.140 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END OAI31M8HM

MACRO OAI31M4HM
    CLASS CORE ;
    FOREIGN OAI31M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER ME1  ;
        ANTENNAGATEAREA 0.288  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.733  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.020 3.500 1.220 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.000 1.020 3.760 1.220 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER ME1  ;
        ANTENNAGATEAREA 0.288  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.661  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.020 1.900 1.220 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.490 1.020 2.210 1.220 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.342  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.860 1.500 5.060 2.020 ;
        RECT  3.820 1.500 5.060 1.740 ;
        RECT  3.820 1.500 4.020 2.020 ;
        RECT  2.640 1.500 5.060 1.660 ;
        RECT  0.100 0.700 3.540 0.860 ;
        RECT  3.260 0.620 3.540 0.860 ;
        RECT  2.640 0.700 2.840 1.660 ;
        RECT  2.440 0.700 2.840 1.160 ;
        RECT  2.180 0.620 2.460 0.860 ;
        RECT  1.140 0.620 1.420 0.860 ;
        RECT  0.100 0.620 0.380 0.860 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER ME1  ;
        ANTENNAGATEAREA 0.288  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.715  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.020 0.700 1.220 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.270 1.020 1.020 1.220 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.216  LAYER ME1  ;
        ANTENNAGATEAREA 0.216  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.600  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.020 4.700 1.220 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  4.120 1.020 4.980 1.240 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.300 -0.140 4.580 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.460 2.460 1.660 ;
        RECT  0.100 1.460 0.380 2.080 ;
        RECT  1.180 1.460 1.380 2.080 ;
        RECT  1.620 1.900 3.580 2.060 ;
        RECT  0.620 0.300 4.020 0.460 ;
        RECT  0.620 0.300 0.900 0.540 ;
        RECT  1.660 0.300 1.940 0.540 ;
        RECT  2.740 0.300 3.020 0.540 ;
        RECT  3.820 0.300 4.020 0.860 ;
        RECT  4.860 0.480 5.060 0.860 ;
        RECT  3.820 0.700 5.060 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OAI31M4HM

MACRO OAI31M2HM
    CLASS CORE ;
    FOREIGN OAI31M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.625  LAYER ME1  ;
        ANTENNADIFFAREA 0.625  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.800 1.900 2.000 ;
        LAYER ME2 ;
        RECT  1.640 1.800 1.960 2.000 ;
        RECT  1.700 1.240 1.900 2.000 ;
        LAYER ME1 ;
        RECT  0.540 1.800 2.090 2.040 ;
        RECT  0.100 0.700 1.510 0.860 ;
        RECT  1.230 0.620 1.510 0.860 ;
        RECT  0.540 0.700 0.740 2.040 ;
        RECT  0.100 0.320 0.380 0.860 ;
        END
    END Z
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.560  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.300 1.500 1.500 ;
        LAYER ME2 ;
        RECT  1.300 0.800 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.020 1.680 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.330 1.640 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.130 1.200 2.700 1.560 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.310 1.840 2.590 2.540 ;
        RECT  0.100 1.840 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.310 -0.140 2.590 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.670 0.300 2.070 0.460 ;
        RECT  0.670 0.300 0.950 0.540 ;
        RECT  1.790 0.300 2.070 0.650 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI31M2HM

MACRO OAI31M1HM
    CLASS CORE ;
    FOREIGN OAI31M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.516  LAYER ME1  ;
        ANTENNADIFFAREA 0.516  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.800 1.900 2.000 ;
        LAYER ME2 ;
        RECT  1.640 1.800 1.960 2.000 ;
        RECT  1.700 1.240 1.900 2.000 ;
        LAYER ME1 ;
        RECT  0.540 1.800 2.030 2.040 ;
        RECT  0.100 0.700 1.510 0.860 ;
        RECT  1.230 0.620 1.510 0.860 ;
        RECT  0.540 0.700 0.740 2.040 ;
        RECT  0.100 0.320 0.380 0.860 ;
        END
    END Z
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        ANTENNAGATEAREA 0.096  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.983  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.290 1.500 1.490 ;
        LAYER ME2 ;
        RECT  1.300 0.800 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.020 1.680 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.330 1.640 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.130 1.200 2.700 1.560 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.350 1.840 2.630 2.540 ;
        RECT  0.100 1.840 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.310 -0.140 2.590 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.670 0.300 2.070 0.460 ;
        RECT  0.670 0.300 0.950 0.540 ;
        RECT  1.790 0.300 2.070 0.600 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI31M1HM

MACRO OAI31M0HM
    CLASS CORE ;
    FOREIGN OAI31M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.455  LAYER ME1  ;
        ANTENNADIFFAREA 0.455  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.800 1.900 2.000 ;
        LAYER ME2 ;
        RECT  1.640 1.800 1.960 2.000 ;
        RECT  1.700 1.240 1.900 2.000 ;
        LAYER ME1 ;
        RECT  0.540 1.800 2.030 2.040 ;
        RECT  0.100 0.700 1.510 0.860 ;
        RECT  1.230 0.620 1.510 0.860 ;
        RECT  0.540 0.700 0.740 2.040 ;
        RECT  0.100 0.380 0.380 0.860 ;
        END
    END Z
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.040  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.300 1.500 1.500 ;
        LAYER ME2 ;
        RECT  1.300 0.760 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.020 1.680 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.330 1.640 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.130 1.200 2.700 1.560 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.350 1.840 2.630 2.540 ;
        RECT  0.100 1.840 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.310 -0.140 2.590 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.670 0.300 2.070 0.460 ;
        RECT  0.670 0.300 0.950 0.540 ;
        RECT  1.790 0.300 2.070 0.540 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI31M0HM

MACRO OAI22M8HM
    CLASS CORE ;
    FOREIGN OAI22M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.363  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.500 1.020 6.700 1.220 ;
        LAYER ME2 ;
        RECT  6.500 0.840 6.700 1.560 ;
        LAYER ME1 ;
        RECT  5.510 1.020 6.830 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.616  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.700 1.020 7.900 1.220 ;
        LAYER ME2 ;
        RECT  7.700 0.840 7.900 1.560 ;
        LAYER ME1 ;
        RECT  7.310 1.020 8.920 1.260 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.680 8.900 0.840 ;
        RECT  8.560 0.620 8.900 0.840 ;
        RECT  7.440 0.620 7.760 0.840 ;
        RECT  2.660 1.580 6.700 1.740 ;
        RECT  6.370 0.620 6.680 0.840 ;
        RECT  4.900 0.620 5.560 0.840 ;
        RECT  4.900 0.620 5.100 1.740 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.570  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.020 3.500 1.220 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.620 1.020 4.100 1.290 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.615  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.540 1.020 2.020 1.340 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.580 1.850 8.860 2.540 ;
        RECT  7.460 1.860 7.740 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.500 2.460 1.660 ;
        RECT  2.240 1.500 2.460 2.060 ;
        RECT  2.240 1.900 4.580 2.060 ;
        RECT  0.100 1.500 0.380 2.100 ;
        RECT  1.150 1.500 1.420 2.100 ;
        RECT  6.940 1.500 9.380 1.660 ;
        RECT  6.940 1.500 7.220 2.100 ;
        RECT  4.740 1.900 7.220 2.100 ;
        RECT  9.100 1.500 9.380 2.100 ;
        RECT  4.260 0.300 9.380 0.460 ;
        RECT  5.790 0.300 6.130 0.500 ;
        RECT  6.920 0.300 7.250 0.500 ;
        RECT  8.000 0.300 8.320 0.500 ;
        RECT  9.100 0.300 9.380 0.680 ;
        RECT  0.160 0.340 0.320 0.860 ;
        RECT  1.200 0.340 1.360 0.860 ;
        RECT  2.240 0.340 2.400 0.860 ;
        RECT  3.280 0.340 3.440 0.860 ;
        RECT  4.260 0.300 4.540 0.860 ;
        RECT  0.160 0.700 4.540 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
    END
END OAI22M8HM

MACRO OAI22M4HM
    CLASS CORE ;
    FOREIGN OAI22M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.780  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.030 3.500 1.230 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.860 1.030 3.650 1.230 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.672  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 1.020 1.680 1.230 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.390 4.340 1.560 ;
        RECT  3.960 1.070 4.340 1.560 ;
        RECT  2.400 1.070 2.700 1.560 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.400 2.140 1.560 ;
        RECT  1.860 1.070 2.140 1.560 ;
        RECT  0.500 1.070 0.780 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.012  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.760 4.700 1.920 ;
        RECT  4.500 0.700 4.700 1.920 ;
        RECT  2.740 0.700 4.700 0.860 ;
        RECT  3.780 0.620 4.060 0.860 ;
        RECT  2.740 0.620 3.020 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.340 2.080 4.620 2.540 ;
        RECT  2.120 2.080 2.400 2.540 ;
        RECT  0.380 1.780 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  1.700 -0.140 1.980 0.540 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.280 0.300 4.580 0.460 ;
        RECT  3.260 0.300 3.540 0.540 ;
        RECT  4.300 0.300 4.580 0.540 ;
        RECT  0.200 0.460 0.360 0.860 ;
        RECT  1.240 0.460 1.400 0.860 ;
        RECT  2.280 0.300 2.440 0.860 ;
        RECT  0.200 0.700 2.440 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OAI22M4HM

MACRO OAI22M2HM
    CLASS CORE ;
    FOREIGN OAI22M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.000 1.540 1.600 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 1.060 2.300 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.000 1.100 1.600 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.640 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.578  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.620 2.700 1.900 ;
        RECT  1.700 1.740 2.700 1.900 ;
        RECT  1.620 0.620 2.700 0.780 ;
        RECT  1.040 1.900 1.860 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.020 2.060 2.300 2.540 ;
        RECT  0.180 1.740 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.540 0.460 ;
        RECT  0.140 0.400 0.340 0.840 ;
        RECT  1.180 0.300 1.380 0.840 ;
        RECT  0.140 0.680 1.380 0.840 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI22M2HM

MACRO OAI22M1HM
    CLASS CORE ;
    FOREIGN OAI22M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.000 1.540 1.600 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 1.060 2.300 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.000 1.100 1.600 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.640 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.483  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.620 2.700 1.900 ;
        RECT  1.700 1.740 2.700 1.900 ;
        RECT  1.660 0.620 2.700 0.780 ;
        RECT  1.040 1.900 1.860 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.020 2.060 2.300 2.540 ;
        RECT  0.180 1.740 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.620 0.460 ;
        RECT  0.140 0.300 0.340 0.840 ;
        RECT  1.180 0.300 1.380 0.840 ;
        RECT  0.140 0.680 1.380 0.840 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.480 2.400 ;
        RECT  2.200 1.140 2.800 2.400 ;
        RECT  0.000 1.200 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
        RECT  1.480 0.000 2.200 1.200 ;
    END
END OAI22M1HM

MACRO OAI22M0HM
    CLASS CORE ;
    FOREIGN OAI22M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.000 1.540 1.600 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 1.060 2.300 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.000 1.100 1.600 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.640 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.429  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.620 2.700 1.900 ;
        RECT  1.700 1.740 2.700 1.900 ;
        RECT  1.660 0.620 2.700 0.780 ;
        RECT  1.040 1.900 1.860 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.020 2.060 2.300 2.540 ;
        RECT  0.180 1.840 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.620 0.460 ;
        RECT  0.140 0.300 0.340 0.840 ;
        RECT  1.180 0.300 1.380 0.840 ;
        RECT  0.140 0.680 1.380 0.840 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.480 2.400 ;
        RECT  2.200 1.140 2.800 2.400 ;
        RECT  0.000 1.200 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
        RECT  1.480 0.000 2.200 1.200 ;
    END
END OAI22M0HM

MACRO OAI22B20M8HM
    CLASS CORE ;
    FOREIGN OAI22B20M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.579  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.060 7.100 1.260 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.200 1.100 7.760 1.260 ;
        RECT  6.840 1.060 7.160 1.260 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.032  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.060 5.500 1.260 ;
        LAYER ME2 ;
        RECT  5.300 0.840 5.500 1.560 ;
        LAYER ME1 ;
        RECT  4.900 1.100 5.850 1.260 ;
        RECT  5.240 1.060 5.560 1.260 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.130  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.540 1.430 ;
        RECT  0.100 1.070 0.300 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.910  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.240 0.690 7.640 0.850 ;
        RECT  7.360 0.620 7.640 0.850 ;
        RECT  6.320 0.620 6.600 0.850 ;
        RECT  5.280 1.450 5.560 1.780 ;
        RECT  5.280 0.620 5.560 0.850 ;
        RECT  4.240 1.450 5.560 1.700 ;
        RECT  3.210 1.200 4.560 1.570 ;
        RECT  4.240 0.690 4.560 1.700 ;
        RECT  4.240 0.620 4.520 1.780 ;
        RECT  3.220 1.200 3.420 1.940 ;
        RECT  2.180 1.540 3.420 1.740 ;
        RECT  2.180 1.540 2.380 1.950 ;
        END
    END Z
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.130  LAYER ME1  ;
        ANTENNAGATEAREA 0.130  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.290  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.070 1.100 1.270 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.740 1.070 1.240 1.390 ;
        END
    END NA1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.360 1.900 7.640 2.540 ;
        RECT  6.320 1.900 6.600 2.540 ;
        RECT  2.660 1.900 2.940 2.540 ;
        RECT  1.140 1.900 1.900 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  3.180 -0.140 3.460 0.530 ;
        RECT  2.200 -0.140 2.400 0.590 ;
        RECT  0.140 -0.140 0.340 0.780 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.980 0.500 1.180 0.910 ;
        RECT  0.980 0.750 1.720 0.910 ;
        RECT  1.520 1.170 2.850 1.330 ;
        RECT  1.520 0.750 1.720 1.710 ;
        RECT  0.660 1.550 1.720 1.710 ;
        RECT  0.660 1.550 0.860 2.030 ;
        RECT  5.800 1.540 8.270 1.740 ;
        RECT  3.720 1.870 4.000 2.100 ;
        RECT  4.760 1.860 5.040 2.100 ;
        RECT  5.800 1.540 6.020 2.100 ;
        RECT  3.720 1.940 6.020 2.100 ;
        RECT  8.050 1.450 8.270 2.100 ;
        RECT  3.700 0.300 8.270 0.460 ;
        RECT  1.580 0.370 2.040 0.530 ;
        RECT  4.760 0.300 5.040 0.530 ;
        RECT  5.800 0.300 6.080 0.530 ;
        RECT  6.840 0.300 7.120 0.530 ;
        RECT  7.990 0.300 8.270 0.530 ;
        RECT  1.880 0.370 2.040 1.000 ;
        RECT  2.720 0.370 2.880 1.000 ;
        RECT  3.700 0.300 3.980 1.000 ;
        RECT  1.880 0.810 3.980 1.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END OAI22B20M8HM

MACRO OAI22B20M4HM
    CLASS CORE ;
    FOREIGN OAI22B20M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.744  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.060 3.900 1.260 ;
        LAYER ME2 ;
        RECT  3.700 1.000 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.530 1.060 4.300 1.260 ;
        END
    END B1
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.464  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.080 1.240 1.280 1.440 ;
        LAYER ME2 ;
        RECT  1.080 1.180 1.500 1.620 ;
        LAYER ME1 ;
        RECT  1.020 1.180 1.350 1.720 ;
        END
    END NA1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.140 1.420 4.700 1.580 ;
        RECT  4.500 1.060 4.700 1.580 ;
        RECT  3.140 1.060 3.340 1.580 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.970 0.460 1.640 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.874  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.300 1.760 5.100 1.920 ;
        RECT  4.900 0.700 5.100 1.920 ;
        RECT  3.260 0.700 5.100 0.860 ;
        RECT  4.300 0.620 4.580 0.860 ;
        RECT  3.260 0.620 3.540 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.660 2.080 4.940 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  1.860 1.750 2.060 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.820 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  2.280 -0.140 2.480 0.600 ;
        RECT  0.140 -0.140 0.340 0.770 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.500 1.180 0.900 ;
        RECT  0.660 0.700 1.670 0.900 ;
        RECT  1.510 0.700 1.670 1.400 ;
        RECT  1.510 1.220 2.810 1.400 ;
        RECT  0.660 0.500 0.860 2.090 ;
        RECT  2.800 0.300 5.100 0.460 ;
        RECT  1.660 0.370 2.120 0.540 ;
        RECT  3.780 0.300 4.060 0.540 ;
        RECT  4.820 0.300 5.100 0.540 ;
        RECT  1.960 0.370 2.120 0.920 ;
        RECT  2.800 0.300 2.960 0.920 ;
        RECT  1.960 0.760 2.960 0.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OAI22B20M4HM

MACRO OAI22B20M2HM
    CLASS CORE ;
    FOREIGN OAI22B20M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.379  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.080 1.300 1.280 1.500 ;
        LAYER ME2 ;
        RECT  0.900 1.240 1.280 1.580 ;
        LAYER ME1 ;
        RECT  1.020 1.180 1.340 1.580 ;
        END
    END NA2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 1.060 2.300 1.560 ;
        RECT  1.920 1.060 2.170 1.720 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.060 2.740 1.600 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.220 0.360 1.640 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.540  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.660 3.100 1.920 ;
        RECT  2.420 1.760 3.100 1.920 ;
        RECT  2.220 0.660 3.100 0.820 ;
        RECT  1.820 1.880 2.580 2.040 ;
        RECT  2.220 0.620 2.500 0.820 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.140 -0.140 1.420 0.660 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.740 2.080 3.020 2.540 ;
        RECT  1.300 1.900 1.580 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.140 0.440 0.340 1.020 ;
        RECT  0.140 0.820 1.720 1.020 ;
        RECT  1.520 0.820 1.720 1.380 ;
        RECT  0.660 0.820 0.860 2.060 ;
        RECT  0.660 1.800 0.980 2.060 ;
        RECT  1.660 0.300 3.060 0.460 ;
        RECT  1.660 0.300 1.940 0.500 ;
        RECT  2.780 0.300 3.060 0.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI22B20M2HM

MACRO OAI22B20M1HM
    CLASS CORE ;
    FOREIGN OAI22B20M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.379  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.080 1.300 1.280 1.500 ;
        LAYER ME2 ;
        RECT  0.900 1.240 1.280 1.580 ;
        LAYER ME1 ;
        RECT  1.020 1.180 1.340 1.580 ;
        END
    END NA2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 1.140 2.300 1.560 ;
        RECT  1.920 1.140 2.170 1.720 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.140 2.740 1.600 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.220 0.360 1.640 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.362  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.820 3.100 1.920 ;
        RECT  2.420 1.760 3.100 1.920 ;
        RECT  2.220 0.820 3.100 0.980 ;
        RECT  1.820 1.880 2.580 2.040 ;
        RECT  2.220 0.620 2.500 0.980 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.140 -0.140 1.420 0.660 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.740 2.080 3.020 2.540 ;
        RECT  1.340 1.900 1.620 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.320 0.440 0.520 1.020 ;
        RECT  0.320 0.820 1.720 1.020 ;
        RECT  1.520 0.820 1.720 1.380 ;
        RECT  0.660 0.820 0.860 2.060 ;
        RECT  0.660 1.800 0.980 2.060 ;
        RECT  1.660 0.300 3.060 0.460 ;
        RECT  1.660 0.300 1.940 0.660 ;
        RECT  2.780 0.300 3.060 0.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI22B20M1HM

MACRO OAI22B20M0HM
    CLASS CORE ;
    FOREIGN OAI22B20M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.379  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.080 1.300 1.280 1.500 ;
        LAYER ME2 ;
        RECT  0.900 1.240 1.280 1.580 ;
        LAYER ME1 ;
        RECT  1.020 1.180 1.340 1.580 ;
        END
    END NA2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 1.140 2.300 1.560 ;
        RECT  1.920 1.140 2.170 1.720 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.140 2.740 1.600 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.220 0.360 1.640 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.325  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.820 3.100 1.920 ;
        RECT  2.420 1.760 3.100 1.920 ;
        RECT  2.220 0.820 3.100 0.980 ;
        RECT  1.820 1.900 2.580 2.060 ;
        RECT  2.220 0.620 2.500 0.980 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.140 -0.140 1.420 0.660 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 2.080 3.100 2.540 ;
        RECT  1.340 1.900 1.620 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.320 0.440 0.520 1.020 ;
        RECT  0.320 0.820 1.720 1.020 ;
        RECT  1.520 0.820 1.720 1.380 ;
        RECT  0.660 0.820 0.860 2.060 ;
        RECT  0.660 1.800 0.980 2.060 ;
        RECT  1.660 0.300 3.060 0.460 ;
        RECT  1.660 0.300 1.940 0.660 ;
        RECT  2.780 0.300 3.060 0.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI22B20M0HM

MACRO OAI22B10M8HM
    CLASS CORE ;
    FOREIGN OAI22B10M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.615  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 0.980 7.100 1.180 ;
        LAYER ME2 ;
        RECT  6.900 0.920 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.240 0.980 7.840 1.140 ;
        RECT  6.840 0.980 7.160 1.180 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.310  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.010 4.700 1.210 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  3.680 1.010 4.940 1.170 ;
        RECT  4.440 1.010 4.760 1.210 ;
        END
    END A1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.998  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.500 7.740 1.660 ;
        RECT  5.300 0.690 5.500 1.660 ;
        RECT  1.620 0.690 5.500 0.850 ;
        RECT  4.860 0.620 5.140 0.850 ;
        RECT  3.820 0.620 4.100 0.850 ;
        RECT  2.660 0.620 2.940 0.850 ;
        RECT  1.620 0.620 1.900 0.850 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.615  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.900 0.980 9.100 1.180 ;
        LAYER ME2 ;
        RECT  8.900 0.920 9.100 1.560 ;
        LAYER ME1 ;
        RECT  8.320 0.980 9.920 1.140 ;
        RECT  8.840 0.980 9.160 1.180 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.726  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.160 1.070 0.360 1.270 ;
        LAYER ME2 ;
        RECT  0.100 0.820 0.360 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.010 0.580 1.310 ;
        END
    END NA2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.500 1.900 9.780 2.540 ;
        RECT  8.460 1.900 8.740 2.540 ;
        RECT  2.660 1.900 2.940 2.540 ;
        RECT  1.620 1.900 1.900 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.500 -0.140 9.780 0.500 ;
        RECT  8.460 -0.140 8.740 0.500 ;
        RECT  7.420 -0.140 7.700 0.500 ;
        RECT  6.380 -0.140 6.660 0.500 ;
        RECT  0.140 -0.140 0.340 0.740 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.510 0.940 0.710 ;
        RECT  0.740 1.010 3.080 1.170 ;
        RECT  0.740 0.510 0.940 2.080 ;
        RECT  0.620 1.520 0.940 2.080 ;
        RECT  1.100 1.500 3.580 1.700 ;
        RECT  3.360 1.500 3.580 2.100 ;
        RECT  1.100 1.500 1.320 2.080 ;
        RECT  2.180 1.500 2.380 2.080 ;
        RECT  3.360 1.900 5.660 2.100 ;
        RECT  1.140 0.300 6.080 0.460 ;
        RECT  2.140 0.300 2.420 0.530 ;
        RECT  3.240 0.300 3.520 0.530 ;
        RECT  4.340 0.300 4.620 0.530 ;
        RECT  5.920 0.300 6.080 0.820 ;
        RECT  6.960 0.400 7.120 0.820 ;
        RECT  8.000 0.400 8.160 0.820 ;
        RECT  9.040 0.400 9.200 0.820 ;
        RECT  1.140 0.300 1.340 0.750 ;
        RECT  10.080 0.400 10.240 0.820 ;
        RECT  5.920 0.660 10.240 0.820 ;
        RECT  7.940 1.500 10.300 1.700 ;
        RECT  9.020 1.500 9.220 2.080 ;
        RECT  10.020 1.500 10.300 2.080 ;
        RECT  7.940 1.500 8.230 2.100 ;
        RECT  5.860 1.900 8.230 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.140 ;
    END
END OAI22B10M8HM

MACRO OAI22B10M4HM
    CLASS CORE ;
    FOREIGN OAI22B10M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.546  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.010 2.300 1.210 ;
        LAYER ME2 ;
        RECT  2.100 0.670 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.960 1.010 2.600 1.230 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.230 0.900 4.900 1.160 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 1.380 5.580 1.540 ;
        RECT  5.080 0.900 5.580 1.540 ;
        RECT  3.700 1.060 3.980 1.540 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.140 0.500 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.031  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.700 4.760 1.900 ;
        RECT  2.100 1.760 3.520 1.920 ;
        RECT  3.260 0.780 3.420 1.920 ;
        RECT  2.830 0.780 3.420 0.940 ;
        RECT  1.620 0.690 3.060 0.850 ;
        RECT  2.780 0.620 3.060 0.850 ;
        RECT  1.620 0.620 1.900 0.850 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.380 1.910 5.660 2.540 ;
        RECT  3.040 2.080 3.720 2.540 ;
        RECT  1.340 1.790 1.540 2.540 ;
        RECT  0.140 1.740 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  4.980 -0.140 5.260 0.320 ;
        RECT  3.860 -0.140 4.140 0.320 ;
        RECT  0.140 -0.140 0.340 0.780 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.820 1.100 3.100 1.300 ;
        RECT  1.460 1.110 1.740 1.580 ;
        RECT  2.820 1.100 2.980 1.580 ;
        RECT  0.680 1.420 2.980 1.580 ;
        RECT  0.680 0.460 0.840 2.050 ;
        RECT  1.140 0.300 3.700 0.460 ;
        RECT  2.160 0.300 2.440 0.530 ;
        RECT  3.240 0.300 3.700 0.530 ;
        RECT  5.510 0.300 5.820 0.650 ;
        RECT  3.540 0.490 5.820 0.650 ;
        RECT  1.140 0.300 1.340 0.770 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END OAI22B10M4HM

MACRO OAI22B10M2HM
    CLASS CORE ;
    FOREIGN OAI22B10M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.060 1.540 1.670 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.060 1.100 1.670 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.700 1.560 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.100 1.180 3.500 1.580 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.566  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 0.620 1.940 0.840 ;
        RECT  1.040 1.840 1.900 2.000 ;
        RECT  1.700 0.620 1.900 2.000 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.260 1.740 3.460 2.540 ;
        RECT  2.060 1.810 2.260 2.540 ;
        RECT  0.180 1.800 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.260 -0.140 3.460 0.800 ;
        RECT  0.620 -0.140 0.900 0.530 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.420 0.460 ;
        RECT  2.220 0.300 2.420 0.680 ;
        RECT  0.140 0.400 0.340 0.850 ;
        RECT  1.180 0.300 1.380 0.850 ;
        RECT  0.140 0.690 1.380 0.850 ;
        RECT  2.060 1.050 2.940 1.330 ;
        RECT  2.740 0.520 2.940 2.010 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI22B10M2HM

MACRO OAI22B10M1HM
    CLASS CORE ;
    FOREIGN OAI22B10M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.110 1.540 1.680 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.110 1.100 1.680 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.130 0.700 1.560 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.100 1.180 3.500 1.580 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.464  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.620 1.980 0.840 ;
        RECT  1.040 1.840 1.900 2.000 ;
        RECT  1.700 0.620 1.900 2.000 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.260 1.780 3.460 2.540 ;
        RECT  2.060 1.740 2.260 2.540 ;
        RECT  0.220 1.740 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.260 -0.140 3.460 0.820 ;
        RECT  0.620 -0.140 0.900 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.680 0.460 ;
        RECT  0.140 0.370 0.340 0.880 ;
        RECT  1.180 0.300 1.380 0.880 ;
        RECT  0.140 0.720 1.380 0.880 ;
        RECT  2.720 0.710 2.940 1.280 ;
        RECT  2.060 1.000 2.940 1.280 ;
        RECT  2.740 0.710 2.940 2.050 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        RECT  3.200 1.140 3.600 2.400 ;
        RECT  0.000 1.290 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  2.400 0.000 3.200 1.290 ;
    END
END OAI22B10M1HM

MACRO OAI22B10M0HM
    CLASS CORE ;
    FOREIGN OAI22B10M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.537  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.180 0.700 1.380 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.720 ;
        LAYER ME1 ;
        RECT  0.100 1.120 0.700 1.440 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.100 1.540 1.740 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.100 1.100 1.740 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.500 1.560 ;
        RECT  3.100 1.040 3.500 1.320 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.620 1.980 0.840 ;
        RECT  1.040 1.930 1.900 2.090 ;
        RECT  1.700 0.620 1.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.260 1.730 3.460 2.540 ;
        RECT  2.060 1.740 2.260 2.540 ;
        RECT  0.220 1.810 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.260 -0.140 3.460 0.840 ;
        RECT  0.620 -0.140 0.900 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.540 0.460 ;
        RECT  2.340 0.300 2.540 0.600 ;
        RECT  0.140 0.400 0.340 0.940 ;
        RECT  1.180 0.300 1.380 0.940 ;
        RECT  0.140 0.780 1.380 0.940 ;
        RECT  2.720 0.800 2.940 1.360 ;
        RECT  2.060 1.080 2.940 1.360 ;
        RECT  2.740 0.800 2.940 2.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.360 2.400 ;
        RECT  0.000 1.380 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  2.360 0.000 3.600 1.380 ;
    END
END OAI22B10M0HM

MACRO OAI222M8HM
    CLASS CORE ;
    FOREIGN OAI222M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 0.909  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.060 8.300 1.260 ;
        LAYER ME2 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  7.980 1.060 8.820 1.260 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.500 1.060 10.700 1.260 ;
        LAYER ME2 ;
        RECT  10.500 0.840 10.700 1.560 ;
        LAYER ME1 ;
        RECT  9.900 1.060 11.380 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.980 1.060 13.900 1.260 ;
        RECT  13.640 0.840 13.900 1.260 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.528  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.300 0.740 13.380 0.900 ;
        RECT  13.100 0.620 13.380 0.900 ;
        RECT  12.060 0.620 12.340 0.900 ;
        RECT  11.020 0.620 11.300 0.900 ;
        RECT  11.060 1.440 11.260 1.720 ;
        RECT  7.460 1.440 11.260 1.600 ;
        RECT  9.980 0.620 10.260 0.900 ;
        RECT  10.020 1.440 10.220 1.720 ;
        RECT  9.300 0.740 9.500 1.600 ;
        RECT  8.500 1.440 8.700 1.720 ;
        RECT  7.460 1.250 7.670 1.600 ;
        RECT  7.460 1.250 7.660 1.720 ;
        RECT  5.330 1.250 7.670 1.410 ;
        RECT  2.740 1.440 5.490 1.600 ;
        RECT  5.330 1.250 5.490 1.600 ;
        RECT  3.780 1.440 3.980 1.720 ;
        RECT  2.740 1.440 2.940 1.720 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 0.804  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.860 1.060 5.060 1.260 ;
        LAYER ME2 ;
        RECT  4.820 0.840 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.450 1.060 5.170 1.260 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.060 3.500 1.260 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.620 1.060 4.100 1.260 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.060 1.500 1.260 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.540 1.060 2.020 1.260 ;
        END
    END C2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.100 1.900 13.380 2.540 ;
        RECT  12.060 1.900 12.340 2.540 ;
        RECT  6.380 1.890 6.660 2.540 ;
        RECT  5.300 2.080 5.580 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  4.260 -0.140 4.540 0.580 ;
        RECT  3.220 -0.140 3.500 0.580 ;
        RECT  2.180 -0.140 2.460 0.580 ;
        RECT  1.140 -0.140 1.420 0.580 ;
        RECT  0.140 -0.140 0.340 0.760 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.540 2.460 1.740 ;
        RECT  2.240 1.540 2.460 2.060 ;
        RECT  4.260 1.810 4.540 2.060 ;
        RECT  2.240 1.900 4.540 2.060 ;
        RECT  0.660 0.480 0.860 0.900 ;
        RECT  1.700 0.480 1.900 0.900 ;
        RECT  2.740 0.480 2.940 0.900 ;
        RECT  3.780 0.480 3.980 0.900 ;
        RECT  5.340 0.620 5.620 0.900 ;
        RECT  6.380 0.620 6.660 0.900 ;
        RECT  7.420 0.620 7.700 0.900 ;
        RECT  8.460 0.620 8.740 0.900 ;
        RECT  0.660 0.740 8.740 0.900 ;
        RECT  5.710 1.570 7.140 1.730 ;
        RECT  5.710 1.570 5.870 1.920 ;
        RECT  4.700 1.760 5.870 1.920 ;
        RECT  6.940 1.570 7.140 2.100 ;
        RECT  7.940 1.820 8.220 2.100 ;
        RECT  8.980 1.820 9.260 2.100 ;
        RECT  6.940 1.940 9.260 2.100 ;
        RECT  11.570 1.540 13.900 1.740 ;
        RECT  9.460 1.820 9.740 2.100 ;
        RECT  10.500 1.820 10.780 2.100 ;
        RECT  11.570 1.540 11.790 2.100 ;
        RECT  9.460 1.940 11.790 2.100 ;
        RECT  4.820 0.300 13.900 0.460 ;
        RECT  4.820 0.300 5.100 0.580 ;
        RECT  5.860 0.300 6.140 0.580 ;
        RECT  6.900 0.300 7.180 0.580 ;
        RECT  7.940 0.300 8.220 0.580 ;
        RECT  8.980 0.300 9.260 0.580 ;
        RECT  9.460 0.300 9.740 0.580 ;
        RECT  10.500 0.300 10.780 0.580 ;
        RECT  11.540 0.300 11.820 0.580 ;
        RECT  12.580 0.300 12.860 0.580 ;
        RECT  13.620 0.300 13.900 0.580 ;
        LAYER VTPH ;
        RECT  0.000 1.140 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.140 ;
    END
END OAI222M8HM

MACRO OAI222M4HM
    CLASS CORE ;
    FOREIGN OAI222M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.000 5.900 1.200 ;
        LAYER ME2 ;
        RECT  5.700 0.840 5.900 1.560 ;
        LAYER ME1 ;
        RECT  5.600 1.000 6.240 1.200 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.000 3.900 1.200 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.520 1.000 4.160 1.200 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.368  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.500 1.060 6.700 1.260 ;
        LAYER ME2 ;
        RECT  6.500 0.840 6.700 1.560 ;
        LAYER ME1 ;
        RECT  5.120 1.360 6.740 1.520 ;
        RECT  6.460 1.000 6.740 1.520 ;
        RECT  5.120 1.000 5.400 1.520 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.020 1.360 4.760 1.520 ;
        RECT  4.400 1.000 4.760 1.520 ;
        RECT  3.020 1.000 3.300 1.520 ;
        END
    END B2
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.360 2.100 1.520 ;
        RECT  1.820 1.000 2.100 1.520 ;
        RECT  0.440 1.000 0.740 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.264  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.100 1.680 7.100 1.840 ;
        RECT  6.900 0.660 7.100 1.840 ;
        RECT  5.260 0.660 7.100 0.820 ;
        RECT  6.300 0.620 6.580 0.820 ;
        RECT  5.260 0.620 5.540 0.820 ;
        END
    END Z
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.000 1.500 1.200 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 1.000 1.600 1.200 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.660 2.080 6.940 2.540 ;
        RECT  4.740 2.080 5.020 2.540 ;
        RECT  2.820 2.080 3.100 2.540 ;
        RECT  2.020 2.080 2.300 2.540 ;
        RECT  0.340 1.780 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.750 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.540 0.900 0.820 ;
        RECT  1.660 0.540 1.940 0.820 ;
        RECT  3.180 0.620 3.460 0.820 ;
        RECT  4.220 0.620 4.500 0.820 ;
        RECT  0.620 0.660 4.500 0.820 ;
        RECT  2.660 0.300 7.100 0.460 ;
        RECT  2.660 0.300 2.940 0.500 ;
        RECT  3.700 0.300 3.980 0.500 ;
        RECT  4.740 0.300 5.020 0.500 ;
        RECT  5.780 0.300 6.060 0.500 ;
        RECT  6.820 0.300 7.100 0.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END OAI222M4HM

MACRO OAI222M2HM
    CLASS CORE ;
    FOREIGN OAI222M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.866  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.000 3.900 1.200 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.360 1.000 3.960 1.220 ;
        END
    END A2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.726  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.010 1.100 1.210 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.000 1.400 1.220 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.726  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.010 1.900 1.210 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.640 1.000 2.200 1.220 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 1.000 3.160 1.320 ;
        RECT  2.880 1.000 3.140 1.780 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.000 2.700 1.780 ;
        END
    END B1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.680 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.500 4.300 1.700 ;
        RECT  4.120 0.660 4.300 1.700 ;
        RECT  3.180 0.660 4.300 0.820 ;
        RECT  2.080 1.940 3.500 2.100 ;
        RECT  3.300 1.500 3.500 2.100 ;
        RECT  3.180 0.620 3.460 0.820 ;
        RECT  2.080 1.540 2.240 2.100 ;
        RECT  1.140 1.540 2.240 1.740 ;
        RECT  1.140 1.540 1.360 1.980 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.660 1.860 3.860 2.540 ;
        RECT  1.720 1.900 1.920 2.540 ;
        RECT  0.300 1.900 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.760 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.540 0.900 0.820 ;
        RECT  2.140 0.620 2.420 0.820 ;
        RECT  0.620 0.660 2.420 0.820 ;
        RECT  1.620 0.300 3.980 0.460 ;
        RECT  1.620 0.300 1.900 0.500 ;
        RECT  2.660 0.300 2.940 0.500 ;
        RECT  3.700 0.300 3.980 0.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OAI222M2HM

MACRO OAI222M1HM
    CLASS CORE ;
    FOREIGN OAI222M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.080 3.900 1.280 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.300 1.060 3.960 1.280 ;
        END
    END A2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.080 1.100 1.280 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.060 1.400 1.280 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.080 1.900 1.280 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.640 1.060 2.200 1.280 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.880 3.100 1.780 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.060 2.700 1.780 ;
        RECT  2.400 1.060 2.700 1.280 ;
        END
    END B1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.680 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.660  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.580 4.300 1.740 ;
        RECT  4.120 0.740 4.300 1.740 ;
        RECT  3.300 0.740 4.300 0.900 ;
        RECT  3.300 0.620 3.580 0.900 ;
        RECT  2.080 1.940 3.500 2.100 ;
        RECT  3.300 1.580 3.500 2.100 ;
        RECT  2.080 1.580 2.280 2.100 ;
        RECT  1.180 1.580 2.280 1.740 ;
        RECT  1.180 1.580 1.380 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.660 1.900 3.860 2.540 ;
        RECT  1.720 1.900 1.920 2.540 ;
        RECT  0.340 1.740 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.580 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.400 0.860 0.900 ;
        RECT  2.180 0.620 2.460 0.900 ;
        RECT  0.660 0.740 2.460 0.900 ;
        RECT  1.620 0.300 4.140 0.460 ;
        RECT  1.620 0.300 1.900 0.580 ;
        RECT  3.860 0.300 4.140 0.580 ;
        RECT  2.780 0.300 2.980 0.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OAI222M1HM

MACRO OAI222M0HM
    CLASS CORE ;
    FOREIGN OAI222M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        ANTENNAGATEAREA 0.082  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.608  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.070 3.900 1.270 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.300 1.060 3.960 1.280 ;
        END
    END A2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        ANTENNAGATEAREA 0.082  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.971  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.070 1.100 1.270 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.060 1.400 1.280 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        ANTENNAGATEAREA 0.082  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.971  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.070 1.900 1.270 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.640 1.060 2.200 1.280 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 1.000 3.100 1.780 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.060 2.700 1.780 ;
        END
    END B1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.680 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.541  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.580 4.300 1.740 ;
        RECT  4.120 0.740 4.300 1.740 ;
        RECT  3.300 0.740 4.300 0.900 ;
        RECT  3.300 0.620 3.580 0.900 ;
        RECT  2.080 1.940 3.500 2.100 ;
        RECT  3.300 1.580 3.500 2.100 ;
        RECT  2.080 1.580 2.240 2.100 ;
        RECT  1.180 1.580 2.240 1.740 ;
        RECT  1.180 1.580 1.380 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.660 1.900 3.860 2.540 ;
        RECT  1.720 1.900 1.920 2.540 ;
        RECT  0.340 1.790 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.580 ;
        RECT  0.140 -0.140 0.340 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.360 0.860 0.900 ;
        RECT  2.180 0.620 2.460 0.900 ;
        RECT  0.660 0.740 2.460 0.900 ;
        RECT  1.620 0.300 4.140 0.460 ;
        RECT  1.620 0.300 1.900 0.580 ;
        RECT  3.860 0.300 4.140 0.580 ;
        RECT  2.780 0.300 2.980 0.640 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OAI222M0HM

MACRO OAI221M8HM
    CLASS CORE ;
    FOREIGN OAI221M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.060 8.300 1.260 ;
        LAYER ME2 ;
        RECT  8.100 0.830 8.300 1.560 ;
        LAYER ME1 ;
        RECT  7.380 1.060 8.860 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.100 1.060 10.300 1.260 ;
        LAYER ME2 ;
        RECT  10.100 0.830 10.300 1.560 ;
        LAYER ME1 ;
        RECT  9.460 1.060 10.940 1.260 ;
        END
    END A2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 2.020 1.260 ;
        RECT  0.100 1.060 0.360 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.438  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.900 0.740 10.860 0.900 ;
        RECT  10.580 0.620 10.860 0.900 ;
        RECT  9.540 0.620 9.820 0.900 ;
        RECT  6.900 1.500 8.820 1.660 ;
        RECT  8.500 0.620 8.780 0.900 ;
        RECT  7.460 0.620 7.740 0.900 ;
        RECT  4.860 1.540 7.100 1.700 ;
        RECT  6.900 0.740 7.100 1.700 ;
        RECT  0.660 1.440 5.220 1.600 ;
        RECT  1.700 1.440 1.900 1.940 ;
        RECT  0.660 1.440 0.860 1.940 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.060 5.900 1.260 ;
        LAYER ME2 ;
        RECT  5.700 0.830 5.900 1.560 ;
        LAYER ME1 ;
        RECT  4.820 1.060 6.300 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.782  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.060 3.500 1.260 ;
        LAYER ME2 ;
        RECT  3.300 0.830 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.480 1.060 4.320 1.260 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.580 1.900 10.860 2.540 ;
        RECT  9.540 1.900 9.820 2.540 ;
        RECT  3.820 2.080 4.100 2.540 ;
        RECT  2.700 2.080 2.980 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  1.660 -0.140 1.940 0.580 ;
        RECT  0.620 -0.140 0.900 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.100 1.760 4.620 1.920 ;
        RECT  4.420 1.880 6.740 2.080 ;
        RECT  0.140 0.480 0.340 0.900 ;
        RECT  1.180 0.480 1.380 0.900 ;
        RECT  2.280 0.480 2.480 0.900 ;
        RECT  3.340 0.620 3.620 0.900 ;
        RECT  4.380 0.620 4.660 0.900 ;
        RECT  5.420 0.620 5.700 0.900 ;
        RECT  6.460 0.620 6.740 0.900 ;
        RECT  0.140 0.740 6.740 0.900 ;
        RECT  2.820 0.300 11.380 0.460 ;
        RECT  2.820 0.300 3.100 0.580 ;
        RECT  3.860 0.300 4.140 0.580 ;
        RECT  4.900 0.300 5.180 0.580 ;
        RECT  5.940 0.300 6.220 0.580 ;
        RECT  6.940 0.300 7.220 0.580 ;
        RECT  7.980 0.300 8.260 0.580 ;
        RECT  9.020 0.300 9.300 0.580 ;
        RECT  10.060 0.300 10.340 0.580 ;
        RECT  11.100 0.300 11.380 0.580 ;
        RECT  9.060 1.540 11.420 1.740 ;
        RECT  9.060 1.540 9.260 2.060 ;
        RECT  6.900 1.900 9.260 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.140 ;
    END
END OAI221M8HM

MACRO OAI221M4HM
    CLASS CORE ;
    FOREIGN OAI221M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.608  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.060 5.100 1.260 ;
        LAYER ME2 ;
        RECT  4.900 0.840 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.760 1.060 5.480 1.260 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.608  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.060 2.700 1.260 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.200 1.060 2.920 1.260 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.320 1.420 5.900 1.580 ;
        RECT  5.700 1.060 5.900 1.580 ;
        RECT  4.320 1.060 4.520 1.580 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.420 3.340 1.580 ;
        RECT  3.140 1.060 3.340 1.580 ;
        RECT  1.700 1.060 1.940 1.580 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.120 1.360 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.175  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.820 1.740 6.300 1.900 ;
        RECT  6.100 0.740 6.300 1.900 ;
        RECT  4.460 0.740 6.300 0.900 ;
        RECT  5.500 0.620 5.780 0.900 ;
        RECT  4.460 0.620 4.740 0.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.860 2.080 6.140 2.540 ;
        RECT  4.100 2.080 4.380 2.540 ;
        RECT  3.300 2.080 3.580 2.540 ;
        RECT  1.480 2.080 1.760 2.540 ;
        RECT  0.380 1.750 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  0.860 -0.140 1.140 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 0.480 0.580 0.900 ;
        RECT  1.420 0.480 1.620 0.900 ;
        RECT  2.420 0.620 2.700 0.900 ;
        RECT  3.460 0.620 3.740 0.900 ;
        RECT  0.380 0.740 3.740 0.900 ;
        RECT  1.900 0.300 6.300 0.460 ;
        RECT  1.900 0.300 2.180 0.580 ;
        RECT  2.940 0.300 3.220 0.580 ;
        RECT  4.980 0.300 5.260 0.580 ;
        RECT  6.020 0.300 6.300 0.580 ;
        RECT  3.980 0.300 4.180 0.760 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END OAI221M4HM

MACRO OAI221M2HM
    CLASS CORE ;
    FOREIGN OAI221M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.020 3.140 1.600 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.020 2.600 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.100 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.020 1.900 1.560 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.700 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.738  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 0.700 3.500 1.920 ;
        RECT  1.260 1.760 3.500 1.920 ;
        RECT  2.700 0.700 3.500 0.860 ;
        RECT  2.700 0.620 2.980 0.860 ;
        RECT  0.620 1.900 1.420 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  1.580 2.080 2.420 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.480 0.860 0.860 ;
        RECT  1.660 0.620 1.940 0.860 ;
        RECT  0.660 0.700 1.940 0.860 ;
        RECT  1.140 0.300 3.500 0.460 ;
        RECT  1.140 0.300 1.420 0.540 ;
        RECT  3.220 0.300 3.500 0.540 ;
        RECT  2.220 0.300 2.420 0.600 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI221M2HM

MACRO OAI221M1HM
    CLASS CORE ;
    FOREIGN OAI221M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 0.960 0.700 1.560 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.060 3.140 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.060 2.600 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.960 1.100 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.080 1.800 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.579  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 0.740 3.500 1.920 ;
        RECT  1.260 1.760 3.500 1.920 ;
        RECT  2.660 0.740 3.500 0.900 ;
        RECT  2.660 0.620 2.940 0.900 ;
        RECT  0.620 1.900 1.420 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  1.580 2.080 2.420 2.540 ;
        RECT  0.140 1.820 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.300 3.500 0.460 ;
        RECT  3.220 0.300 3.500 0.580 ;
        RECT  2.140 0.300 2.340 0.670 ;
        RECT  1.140 0.300 1.420 0.800 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.460 2.400 ;
        RECT  2.200 1.140 3.600 2.400 ;
        RECT  0.000 1.280 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  0.460 0.000 2.200 1.280 ;
    END
END OAI221M1HM

MACRO OAI221M0HM
    CLASS CORE ;
    FOREIGN OAI221M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.960 0.700 1.560 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.060 3.140 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.060 2.600 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 1.020 1.100 1.780 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.060 1.900 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.760 3.500 1.920 ;
        RECT  3.300 0.740 3.500 1.920 ;
        RECT  2.660 0.740 3.500 0.900 ;
        RECT  2.660 0.620 2.940 0.900 ;
        RECT  0.650 1.940 1.420 2.100 ;
        RECT  1.260 1.760 1.420 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.140 2.080 2.420 2.540 ;
        RECT  1.610 2.080 1.890 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  0.140 -0.140 0.340 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.300 3.500 0.460 ;
        RECT  3.220 0.300 3.500 0.580 ;
        RECT  2.140 0.300 2.340 0.650 ;
        RECT  1.140 0.300 1.420 0.800 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.460 2.400 ;
        RECT  2.200 1.140 3.600 2.400 ;
        RECT  0.000 1.230 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  0.460 0.000 2.200 1.230 ;
    END
END OAI221M0HM

MACRO OAI21M8HM
    CLASS CORE ;
    FOREIGN OAI21M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.473  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 1.540 1.270 ;
        RECT  0.100 1.070 0.360 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.820 1.540 4.100 1.780 ;
        RECT  0.740 1.540 4.100 1.700 ;
        RECT  2.780 1.540 3.060 1.780 ;
        RECT  1.780 1.540 2.020 1.940 ;
        RECT  0.700 0.750 2.020 0.910 ;
        RECT  1.740 0.620 2.020 0.910 ;
        RECT  1.700 0.750 1.900 1.700 ;
        RECT  0.700 0.620 0.980 0.910 ;
        RECT  0.740 1.540 0.940 1.950 ;
        END
    END Z
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.435  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.860 1.040 4.260 1.240 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.507  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.040 5.500 1.240 ;
        LAYER ME2 ;
        RECT  5.300 0.840 5.500 1.560 ;
        LAYER ME1 ;
        RECT  4.780 1.040 6.260 1.240 ;
        END
    END A2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.900 1.900 6.180 2.540 ;
        RECT  4.860 1.900 5.140 2.540 ;
        RECT  1.220 1.900 1.500 2.540 ;
        RECT  0.180 1.900 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.900 -0.140 6.180 0.500 ;
        RECT  4.860 -0.140 5.140 0.500 ;
        RECT  3.820 -0.140 4.100 0.500 ;
        RECT  2.780 -0.140 3.060 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.340 1.540 6.700 1.740 ;
        RECT  2.260 1.900 2.540 2.100 ;
        RECT  3.300 1.900 3.580 2.100 ;
        RECT  5.420 1.540 5.620 1.990 ;
        RECT  6.480 1.540 6.700 1.990 ;
        RECT  4.340 1.540 4.560 2.100 ;
        RECT  2.260 1.940 4.560 2.100 ;
        RECT  0.180 0.300 2.340 0.460 ;
        RECT  1.220 0.300 1.500 0.590 ;
        RECT  2.180 0.440 2.620 0.600 ;
        RECT  2.460 0.440 2.620 0.880 ;
        RECT  3.300 0.620 3.580 0.880 ;
        RECT  4.340 0.620 4.620 0.880 ;
        RECT  5.380 0.620 5.660 0.880 ;
        RECT  0.180 0.300 0.460 0.780 ;
        RECT  6.420 0.490 6.700 0.880 ;
        RECT  2.460 0.720 6.700 0.880 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END OAI21M8HM

MACRO OAI21M6HM
    CLASS CORE ;
    FOREIGN OAI21M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.433  LAYER ME1  ;
        ANTENNAGATEAREA 0.433  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.080  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.000 2.300 1.200 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.040 1.000 2.740 1.200 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.433  LAYER ME1  ;
        ANTENNAGATEAREA 0.433  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.536  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 0.980 1.100 1.180 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.520 0.980 1.600 1.180 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.425  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.300 1.480 4.700 2.020 ;
        RECT  2.220 1.480 4.700 1.640 ;
        RECT  3.260 1.480 3.540 2.020 ;
        RECT  2.900 0.620 3.100 1.640 ;
        RECT  0.660 0.660 3.100 0.820 ;
        RECT  2.740 0.620 3.100 0.820 ;
        RECT  2.220 1.480 2.500 1.710 ;
        RECT  1.700 0.620 1.980 0.820 ;
        RECT  0.660 0.620 0.940 0.820 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.352  LAYER ME1  ;
        ANTENNAGATEAREA 0.352  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.011  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.000 3.900 1.200 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.600 1.000 4.760 1.200 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  3.780 1.900 4.060 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.140 1.540 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.860 -0.140 5.060 0.840 ;
        RECT  3.780 -0.140 4.060 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.540 1.980 1.740 ;
        RECT  1.760 1.540 1.980 2.100 ;
        RECT  0.660 1.540 0.880 2.100 ;
        RECT  2.740 1.840 3.020 2.100 ;
        RECT  1.760 1.940 3.020 2.100 ;
        RECT  0.140 0.300 3.480 0.460 ;
        RECT  1.180 0.300 1.460 0.500 ;
        RECT  2.220 0.300 2.500 0.500 ;
        RECT  3.320 0.300 3.480 0.820 ;
        RECT  0.140 0.300 0.420 0.780 ;
        RECT  4.300 0.470 4.580 0.820 ;
        RECT  3.320 0.660 4.580 0.820 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OAI21M6HM

MACRO OAI21M4HM
    CLASS CORE ;
    FOREIGN OAI21M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.528  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.080 2.300 1.280 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.000 1.070 2.640 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 1.440 3.140 1.600 ;
        RECT  2.860 1.070 3.140 1.600 ;
        RECT  1.500 1.070 1.780 1.600 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.070 1.080 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.877  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.580 1.760 3.500 1.920 ;
        RECT  3.300 0.750 3.500 1.920 ;
        RECT  1.660 0.750 3.500 0.910 ;
        RECT  2.700 0.620 2.980 0.910 ;
        RECT  1.660 0.620 1.940 0.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.060 2.080 3.340 2.540 ;
        RECT  1.240 2.080 1.520 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  0.620 -0.140 0.900 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 0.300 3.500 0.460 ;
        RECT  2.180 0.300 2.460 0.590 ;
        RECT  3.220 0.300 3.500 0.590 ;
        RECT  0.160 0.460 0.320 0.910 ;
        RECT  1.200 0.300 1.360 0.910 ;
        RECT  0.160 0.750 1.360 0.910 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI21M4HM

MACRO OAI21M3HM
    CLASS CORE ;
    FOREIGN OAI21M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.217  LAYER ME1  ;
        ANTENNAGATEAREA 0.217  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.011  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 0.980 1.100 1.180 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.820 0.980 1.460 1.180 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 1.440 1.940 1.600 ;
        RECT  1.660 1.000 1.940 1.600 ;
        RECT  0.340 1.170 0.500 1.600 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.000 2.700 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.765  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.960 1.760 3.100 1.920 ;
        RECT  2.900 0.660 3.100 1.920 ;
        RECT  0.320 0.660 3.100 0.820 ;
        RECT  1.440 0.620 1.720 0.820 ;
        RECT  0.320 0.340 0.600 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.880 2.080 2.160 2.540 ;
        RECT  0.140 1.830 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.480 -0.140 2.760 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.920 0.300 2.240 0.460 ;
        RECT  0.920 0.300 1.200 0.500 ;
        RECT  1.960 0.300 2.240 0.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI21M3HM

MACRO OAI21M2HM
    CLASS CORE ;
    FOREIGN OAI21M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.114  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.130 1.900 1.330 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.100 1.960 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.100 1.100 1.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.640 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.576  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.540 2.300 1.740 ;
        RECT  2.120 0.780 2.300 1.740 ;
        RECT  0.620 0.780 2.300 0.940 ;
        RECT  1.040 1.900 1.500 2.100 ;
        RECT  1.300 1.540 1.500 2.100 ;
        RECT  0.620 0.620 0.900 0.940 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.660 -0.140 1.940 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.300 1.420 0.460 ;
        RECT  1.140 0.300 1.420 0.590 ;
        RECT  0.160 0.300 0.320 0.810 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END OAI21M2HM

MACRO OAI21M1HM
    CLASS CORE ;
    FOREIGN OAI21M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.903  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.180 1.900 1.380 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.140 1.960 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.140 1.100 1.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.140 0.700 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.464  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.580 2.300 1.740 ;
        RECT  2.120 0.780 2.300 1.740 ;
        RECT  0.660 0.780 2.300 0.980 ;
        RECT  1.000 1.900 1.500 2.100 ;
        RECT  1.300 1.580 1.500 2.100 ;
        RECT  0.660 0.620 0.940 0.980 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.140 1.740 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.740 -0.140 2.020 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.300 1.500 0.460 ;
        RECT  1.220 0.300 1.500 0.620 ;
        RECT  0.160 0.300 0.320 0.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END OAI21M1HM

MACRO OAI21M0HM
    CLASS CORE ;
    FOREIGN OAI21M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.023  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.180 1.900 1.380 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.140 1.960 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.140 1.100 1.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 1.140 0.700 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.406  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.580 2.300 1.740 ;
        RECT  2.120 0.820 2.300 1.740 ;
        RECT  0.660 0.820 2.300 0.980 ;
        RECT  1.000 1.900 1.500 2.100 ;
        RECT  1.300 1.580 1.500 2.100 ;
        RECT  0.660 0.620 0.940 0.980 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.700 1.900 1.980 2.540 ;
        RECT  0.140 1.770 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.740 -0.140 2.020 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.300 1.500 0.460 ;
        RECT  1.220 0.300 1.500 0.660 ;
        RECT  0.160 0.300 0.320 0.760 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END OAI21M0HM

MACRO OAI21B20M8HM
    CLASS CORE ;
    FOREIGN OAI21B20M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.502  LAYER ME1  ;
        ANTENNAGATEAREA 0.502  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.234  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.140 2.300 1.340 ;
        LAYER ME2 ;
        RECT  2.100 0.930 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.760 1.320 4.320 1.480 ;
        RECT  4.040 1.120 4.320 1.480 ;
        RECT  1.760 1.120 2.400 1.480 ;
        END
    END B
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.130  LAYER ME1  ;
        ANTENNAGATEAREA 0.130  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.210  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.070 1.100 1.270 ;
        LAYER ME2 ;
        RECT  0.900 0.930 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.780 0.980 1.180 1.380 ;
        END
    END NA2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.130  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.500 1.340 ;
        RECT  0.100 1.020 0.360 1.560 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.224  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 1.640 5.100 1.800 ;
        RECT  4.940 0.480 5.100 1.800 ;
        RECT  1.900 0.480 5.100 0.640 ;
        RECT  4.100 1.640 4.360 1.960 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.780 1.960 5.060 2.540 ;
        RECT  3.660 1.960 3.940 2.540 ;
        RECT  2.500 1.960 2.780 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.780 -0.140 5.060 0.320 ;
        RECT  3.020 -0.140 3.300 0.320 ;
        RECT  0.940 -0.140 1.220 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.470 0.380 0.820 ;
        RECT  0.100 0.660 1.500 0.820 ;
        RECT  1.340 0.800 4.780 0.960 ;
        RECT  2.800 0.800 3.520 1.160 ;
        RECT  4.620 0.800 4.780 1.260 ;
        RECT  1.340 0.660 1.500 1.740 ;
        RECT  0.680 1.580 1.500 1.740 ;
        RECT  0.680 1.580 0.840 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OAI21B20M8HM

MACRO OAI21B20M4HM
    CLASS CORE ;
    FOREIGN OAI21B20M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.251  LAYER ME1  ;
        ANTENNAGATEAREA 0.251  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.576  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.060 2.300 1.260 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.900 0.980 2.300 1.340 ;
        END
    END B
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.647  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 0.980 1.100 1.180 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.860 0.920 1.180 1.340 ;
        END
    END NA2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 0.700 1.300 ;
        RECT  0.100 0.980 0.300 1.560 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.612  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.720 1.580 3.500 1.740 ;
        RECT  3.300 0.720 3.500 1.740 ;
        RECT  2.780 0.720 3.500 0.880 ;
        RECT  2.740 1.580 2.940 2.010 ;
        RECT  2.780 0.300 2.940 0.880 ;
        RECT  2.140 0.300 2.940 0.500 ;
        RECT  1.720 1.580 1.920 2.010 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.120 -0.140 3.380 0.560 ;
        RECT  1.240 -0.140 1.520 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.820 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.340 0.310 0.540 0.760 ;
        RECT  0.340 0.560 1.720 0.760 ;
        RECT  1.520 0.660 2.620 0.820 ;
        RECT  2.460 0.660 2.620 1.240 ;
        RECT  2.460 1.040 3.140 1.240 ;
        RECT  1.520 0.560 1.720 1.340 ;
        RECT  1.350 1.140 1.550 1.740 ;
        RECT  0.660 1.580 1.550 1.740 ;
        RECT  0.660 1.580 0.860 2.090 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI21B20M4HM

MACRO OAI21B20M2HM
    CLASS CORE ;
    FOREIGN OAI21B20M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.126  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.000 0.980 1.500 1.300 ;
        END
    END NA2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.730 2.340 1.280 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 0.560 1.560 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.409  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.540 2.700 1.740 ;
        RECT  2.500 0.300 2.700 1.740 ;
        RECT  2.300 0.300 2.700 0.500 ;
        RECT  1.900 1.900 2.260 2.100 ;
        RECT  2.060 1.540 2.260 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.420 1.900 2.700 2.540 ;
        RECT  1.380 1.900 1.660 2.540 ;
        RECT  0.220 1.840 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.400 -0.140 1.680 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.500 0.340 0.780 0.820 ;
        RECT  0.500 0.660 1.860 0.820 ;
        RECT  1.660 0.660 1.860 1.740 ;
        RECT  0.780 1.540 1.860 1.740 ;
        RECT  0.780 1.540 1.060 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI21B20M2HM

MACRO OAI21B20M1HM
    CLASS CORE ;
    FOREIGN OAI21B20M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.023  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.190 1.100 1.390 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.130 1.500 1.410 ;
        END
    END NA2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.088  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.340 1.280 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.130 0.560 1.560 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.301  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.580 2.700 1.740 ;
        RECT  2.500 0.390 2.700 1.740 ;
        RECT  2.340 0.390 2.700 0.590 ;
        RECT  1.900 1.900 2.260 2.100 ;
        RECT  2.060 1.580 2.260 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.420 1.900 2.700 2.540 ;
        RECT  1.380 1.900 1.660 2.540 ;
        RECT  0.220 1.840 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.400 -0.140 1.680 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.540 0.430 0.740 0.970 ;
        RECT  0.540 0.810 1.860 0.970 ;
        RECT  1.700 0.810 1.860 1.740 ;
        RECT  0.780 1.580 1.860 1.740 ;
        RECT  0.780 1.580 1.060 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI21B20M1HM

MACRO OAI21B20M0HM
    CLASS CORE ;
    FOREIGN OAI21B20M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        ANTENNAGATEAREA 0.071  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.023  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.150 1.500 1.350 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.000 1.090 1.500 1.410 ;
        END
    END NA2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.800 2.340 1.410 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.240 1.130 0.700 1.560 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.247  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.580 2.700 1.740 ;
        RECT  2.500 0.350 2.700 1.740 ;
        RECT  2.340 0.350 2.700 0.550 ;
        RECT  1.900 1.900 2.260 2.100 ;
        RECT  2.060 1.580 2.260 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.420 1.900 2.700 2.540 ;
        RECT  1.380 1.900 1.660 2.540 ;
        RECT  0.380 1.840 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.400 -0.140 1.680 0.610 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.540 0.390 0.740 0.930 ;
        RECT  0.540 0.770 1.860 0.930 ;
        RECT  1.660 0.770 1.860 1.740 ;
        RECT  0.860 1.580 1.860 1.740 ;
        RECT  0.860 1.580 1.140 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI21B20M0HM

MACRO OAI21B10M8HM
    CLASS CORE ;
    FOREIGN OAI21B10M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.471  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.000 3.900 1.200 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.520 1.000 4.960 1.200 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.473  LAYER ME1  ;
        ANTENNAGATEAREA 0.473  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.166  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.000 6.300 1.200 ;
        LAYER ME2 ;
        RECT  6.100 0.840 6.300 1.560 ;
        LAYER ME1 ;
        RECT  5.900 1.000 6.640 1.320 ;
        END
    END B
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.290 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.484  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.020 0.680 7.340 0.840 ;
        RECT  7.060 0.620 7.340 0.840 ;
        RECT  6.860 1.490 7.100 1.900 ;
        RECT  6.900 0.680 7.100 1.900 ;
        RECT  5.300 1.490 7.100 1.650 ;
        RECT  6.020 0.620 6.300 0.840 ;
        RECT  5.820 1.490 6.020 1.890 ;
        RECT  3.660 1.500 6.020 1.660 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.340 1.850 7.620 2.540 ;
        RECT  6.300 1.850 6.580 2.540 ;
        RECT  2.660 1.850 2.940 2.540 ;
        RECT  1.620 1.850 1.900 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  4.740 -0.140 5.020 0.500 ;
        RECT  3.700 -0.140 3.980 0.500 ;
        RECT  2.660 -0.140 2.940 0.500 ;
        RECT  1.620 -0.140 1.900 0.500 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.000 3.060 1.160 ;
        RECT  0.660 0.410 0.860 2.080 ;
        RECT  1.100 1.490 3.460 1.690 ;
        RECT  3.240 1.490 3.460 2.100 ;
        RECT  4.220 1.820 4.500 2.100 ;
        RECT  1.100 1.490 1.320 1.940 ;
        RECT  2.180 1.490 2.380 2.020 ;
        RECT  5.260 1.820 5.540 2.100 ;
        RECT  3.240 1.940 5.540 2.100 ;
        RECT  5.520 0.300 7.900 0.460 ;
        RECT  6.540 0.300 6.820 0.500 ;
        RECT  7.620 0.300 7.900 0.500 ;
        RECT  1.100 0.440 1.380 0.820 ;
        RECT  2.140 0.530 2.420 0.820 ;
        RECT  3.180 0.530 3.460 0.820 ;
        RECT  4.220 0.530 4.500 0.820 ;
        RECT  5.520 0.300 5.680 0.820 ;
        RECT  1.100 0.660 5.680 0.820 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END OAI21B10M8HM

MACRO OAI21B10M4HM
    CLASS CORE ;
    FOREIGN OAI21B10M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.510  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.070 3.500 1.270 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.200 1.070 3.840 1.270 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        ANTENNAGATEAREA 0.235  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.034  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.070 1.900 1.270 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.600 1.070 2.320 1.270 ;
        END
    END B
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 1.140 0.700 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.877  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 1.750 4.700 1.910 ;
        RECT  4.500 0.740 4.700 1.910 ;
        RECT  2.860 0.740 4.700 0.900 ;
        RECT  3.900 0.620 4.180 0.900 ;
        RECT  2.860 0.620 3.140 0.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.260 2.070 4.540 2.540 ;
        RECT  2.440 2.070 2.720 2.540 ;
        RECT  1.340 1.780 1.540 2.540 ;
        RECT  0.340 1.720 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  1.820 -0.140 2.100 0.590 ;
        RECT  0.340 -0.140 0.540 0.810 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.700 1.070 2.980 1.590 ;
        RECT  4.100 1.060 4.300 1.590 ;
        RECT  0.880 1.430 4.300 1.590 ;
        RECT  0.880 0.500 1.040 2.020 ;
        RECT  2.400 0.300 4.700 0.460 ;
        RECT  3.380 0.300 3.660 0.580 ;
        RECT  4.420 0.300 4.700 0.580 ;
        RECT  1.360 0.430 1.520 0.910 ;
        RECT  2.400 0.300 2.560 0.910 ;
        RECT  1.360 0.750 2.560 0.910 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OAI21B10M4HM

MACRO OAI21B10M2HM
    CLASS CORE ;
    FOREIGN OAI21B10M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.933  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.120 2.700 1.320 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.400 1.070 2.760 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.070 2.240 1.290 ;
        RECT  1.700 1.070 1.900 1.560 ;
        END
    END A1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.220 0.700 1.540 ;
        RECT  0.100 1.220 0.300 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.440  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.540 3.100 1.740 ;
        RECT  2.920 0.750 3.100 1.740 ;
        RECT  1.620 0.750 3.100 0.910 ;
        RECT  2.100 1.540 2.360 2.020 ;
        RECT  1.620 0.620 1.900 0.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.660 1.900 2.940 2.540 ;
        RECT  1.340 1.680 1.540 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.660 -0.140 2.940 0.590 ;
        RECT  0.140 -0.140 0.340 0.800 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.520 0.860 1.020 ;
        RECT  0.660 0.780 1.100 1.020 ;
        RECT  0.900 1.070 1.540 1.230 ;
        RECT  0.900 0.780 1.100 1.930 ;
        RECT  0.620 1.730 1.100 1.930 ;
        RECT  1.100 0.300 2.420 0.460 ;
        RECT  1.100 0.300 1.380 0.590 ;
        RECT  2.140 0.300 2.420 0.590 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI21B10M2HM

MACRO OAI21B10M1HM
    CLASS CORE ;
    FOREIGN OAI21B10M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.396  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.340 1.100 2.760 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.100 2.180 1.380 ;
        RECT  1.700 1.100 1.900 1.560 ;
        END
    END A1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 1.150 0.700 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.357  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.540 3.100 1.740 ;
        RECT  2.920 0.780 3.100 1.740 ;
        RECT  1.660 0.780 3.100 0.940 ;
        RECT  2.100 1.540 2.360 2.090 ;
        RECT  1.660 0.620 1.940 0.940 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.740 -0.140 3.020 0.620 ;
        RECT  0.140 -0.140 0.340 0.730 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.660 1.900 2.940 2.540 ;
        RECT  1.340 1.740 1.540 2.540 ;
        RECT  0.140 1.720 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.660 0.450 0.860 0.980 ;
        RECT  0.660 0.780 1.100 0.980 ;
        RECT  0.900 1.090 1.540 1.370 ;
        RECT  0.900 0.780 1.100 1.930 ;
        RECT  0.620 1.730 1.100 1.930 ;
        RECT  1.100 0.300 2.500 0.460 ;
        RECT  1.100 0.300 1.380 0.620 ;
        RECT  2.220 0.300 2.500 0.620 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI21B10M1HM

MACRO OAI21B10M0HM
    CLASS CORE ;
    FOREIGN OAI21B10M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.230  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.340 1.100 2.760 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.100 2.180 1.380 ;
        RECT  1.700 1.100 1.900 1.560 ;
        END
    END A1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 1.220 0.760 1.540 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.342  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.540 3.100 1.740 ;
        RECT  2.940 0.780 3.100 1.740 ;
        RECT  1.660 0.780 3.100 0.940 ;
        RECT  2.100 1.540 2.420 2.100 ;
        RECT  1.660 0.620 1.940 0.940 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.740 -0.140 3.020 0.620 ;
        RECT  0.140 -0.140 0.340 0.800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.740 1.900 3.020 2.540 ;
        RECT  1.340 1.770 1.540 2.540 ;
        RECT  0.140 1.700 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.660 0.520 0.860 1.020 ;
        RECT  0.660 0.820 1.100 1.020 ;
        RECT  0.920 1.100 1.540 1.380 ;
        RECT  0.920 0.820 1.100 1.930 ;
        RECT  0.620 1.730 1.100 1.930 ;
        RECT  1.100 0.300 2.500 0.460 ;
        RECT  1.100 0.300 1.380 0.620 ;
        RECT  2.220 0.300 2.500 0.620 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OAI21B10M0HM

MACRO OAI21B01M8HM
    CLASS CORE ;
    FOREIGN OAI21B01M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.938  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.040 5.900 1.240 ;
        LAYER ME2 ;
        RECT  5.700 0.960 5.900 1.560 ;
        LAYER ME1 ;
        RECT  5.540 1.040 7.500 1.240 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.148  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.960 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.120 1.040 4.200 1.240 ;
        END
    END A1
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.800 1.240 ;
        RECT  0.100 0.840 0.300 1.240 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.413  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.380 1.530 4.900 1.690 ;
        RECT  2.440 0.620 2.760 1.690 ;
        RECT  2.420 1.530 2.700 1.770 ;
        RECT  1.380 0.660 2.760 0.820 ;
        RECT  2.420 0.620 2.760 0.820 ;
        RECT  1.380 1.530 1.660 1.830 ;
        RECT  1.380 0.560 1.660 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.660 1.900 6.940 2.540 ;
        RECT  5.620 1.900 5.900 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.660 -0.140 6.940 0.540 ;
        RECT  5.620 -0.140 5.900 0.540 ;
        RECT  4.580 -0.140 4.860 0.540 ;
        RECT  3.500 -0.140 3.780 0.540 ;
        RECT  0.860 -0.140 1.140 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 0.300 0.690 0.580 ;
        RECT  0.530 0.300 0.690 0.820 ;
        RECT  0.530 0.660 1.180 0.820 ;
        RECT  0.980 1.090 2.060 1.290 ;
        RECT  0.980 0.660 1.180 1.700 ;
        RECT  0.340 1.500 1.180 1.700 ;
        RECT  5.140 1.520 7.500 1.720 ;
        RECT  5.140 1.520 5.340 2.060 ;
        RECT  2.980 1.900 5.340 2.060 ;
        RECT  1.880 0.300 3.260 0.460 ;
        RECT  1.880 0.300 2.200 0.500 ;
        RECT  2.900 0.300 3.260 0.500 ;
        RECT  3.100 0.300 3.260 0.860 ;
        RECT  4.060 0.600 4.340 0.860 ;
        RECT  5.100 0.600 5.380 0.860 ;
        RECT  6.140 0.600 6.420 0.860 ;
        RECT  7.220 0.320 7.500 0.860 ;
        RECT  3.100 0.700 7.500 0.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END OAI21B01M8HM

MACRO OAI21B01M4HM
    CLASS CORE ;
    FOREIGN OAI21B01M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.654  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.000 3.900 1.200 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.280 1.000 4.000 1.200 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.700 1.420 4.500 1.580 ;
        RECT  4.220 1.070 4.500 1.580 ;
        RECT  2.700 1.240 3.100 1.580 ;
        RECT  2.700 1.070 2.980 1.580 ;
        END
    END A2
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.140 0.500 1.560 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.674  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 1.740 3.860 1.900 ;
        RECT  1.700 0.620 1.900 1.900 ;
        RECT  1.620 0.620 1.900 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.420 2.060 4.700 2.540 ;
        RECT  2.440 2.060 2.720 2.540 ;
        RECT  1.140 1.800 1.340 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.900 -0.140 4.180 0.500 ;
        RECT  2.860 -0.140 3.140 0.500 ;
        RECT  0.140 -0.140 0.340 0.800 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 1.070 1.540 1.250 ;
        RECT  0.680 0.520 0.880 1.970 ;
        RECT  1.100 0.300 2.380 0.460 ;
        RECT  1.100 0.300 1.380 0.590 ;
        RECT  2.180 0.300 2.380 0.820 ;
        RECT  3.380 0.530 3.660 0.820 ;
        RECT  4.420 0.530 4.700 0.820 ;
        RECT  2.180 0.660 4.700 0.820 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OAI21B01M4HM

MACRO OAI21B01M2HM
    CLASS CORE ;
    FOREIGN OAI21B01M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.060 1.620 1.640 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 1.060 2.320 1.560 ;
        END
    END A2
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.180 0.700 1.560 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.545  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.660 2.700 1.920 ;
        RECT  1.780 1.720 2.700 1.920 ;
        RECT  1.740 0.660 2.700 0.840 ;
        RECT  1.740 0.620 2.140 0.840 ;
        RECT  1.260 1.830 1.920 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.840 ;
        RECT  0.100 0.660 1.100 0.840 ;
        RECT  0.900 0.660 1.100 1.920 ;
        RECT  0.100 1.720 1.100 1.920 ;
        RECT  0.100 1.720 0.380 2.060 ;
        RECT  1.180 0.300 2.620 0.460 ;
        RECT  2.300 0.300 2.620 0.500 ;
        RECT  1.180 0.300 1.540 0.520 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI21B01M2HM

MACRO OAI21B01M1HM
    CLASS CORE ;
    FOREIGN OAI21B01M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.150 1.620 1.640 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.030 1.140 2.320 1.560 ;
        END
    END A2
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.150 0.700 1.560 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.429  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.660 2.700 1.880 ;
        RECT  1.780 1.720 2.700 1.880 ;
        RECT  1.700 0.660 2.700 0.840 ;
        RECT  1.700 0.620 2.140 0.840 ;
        RECT  1.260 1.860 1.940 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.840 ;
        RECT  0.100 0.660 1.090 0.840 ;
        RECT  0.890 0.660 1.090 1.920 ;
        RECT  0.100 1.720 1.090 1.920 ;
        RECT  0.100 1.720 0.380 2.060 ;
        RECT  1.180 0.300 2.620 0.460 ;
        RECT  2.300 0.300 2.620 0.500 ;
        RECT  1.180 0.300 1.540 0.520 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI21B01M1HM

MACRO OAI21B01M0HM
    CLASS CORE ;
    FOREIGN OAI21B01M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.000 1.740 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 1.000 2.340 1.560 ;
        END
    END A2
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.040 0.700 1.560 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.660 2.700 1.920 ;
        RECT  1.780 1.720 2.700 1.920 ;
        RECT  1.780 0.660 2.700 0.840 ;
        RECT  1.780 0.620 2.140 0.840 ;
        RECT  1.260 1.800 1.910 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.840 ;
        RECT  0.100 0.660 1.100 0.840 ;
        RECT  0.860 0.660 1.100 1.920 ;
        RECT  0.100 1.720 1.100 1.920 ;
        RECT  0.100 1.720 0.380 2.060 ;
        RECT  1.180 0.300 2.700 0.460 ;
        RECT  2.380 0.300 2.700 0.500 ;
        RECT  1.180 0.300 1.540 0.520 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OAI21B01M0HM

MACRO OAI211M8HM
    CLASS CORE ;
    FOREIGN OAI211M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.590  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.040 5.500 1.240 ;
        LAYER ME2 ;
        RECT  5.300 0.840 5.500 1.560 ;
        LAYER ME1 ;
        RECT  4.700 0.980 6.220 1.280 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.488  LAYER ME1  ;
        ANTENNAGATEAREA 0.488  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.704  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.040 3.100 1.240 ;
        LAYER ME2 ;
        RECT  2.900 0.840 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.520 0.980 3.720 1.380 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.780 1.000 8.700 1.280 ;
        RECT  8.380 0.660 8.700 1.280 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.253  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 0.660 8.220 0.820 ;
        RECT  7.860 0.620 8.220 0.820 ;
        RECT  6.820 0.620 7.180 0.820 ;
        RECT  5.780 1.540 6.140 1.780 ;
        RECT  5.780 0.620 6.140 0.820 ;
        RECT  0.620 1.540 6.140 1.740 ;
        RECT  4.740 1.540 5.100 1.780 ;
        RECT  4.740 0.620 5.100 0.820 ;
        RECT  4.100 0.660 4.300 1.740 ;
        RECT  3.780 1.540 4.060 2.020 ;
        RECT  2.740 1.540 3.020 2.020 ;
        RECT  1.660 1.540 1.940 2.020 ;
        RECT  0.620 1.540 0.900 1.940 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.488  LAYER ME1  ;
        ANTENNAGATEAREA 0.488  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.554  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.040 1.100 1.240 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.440 1.000 1.600 1.300 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  3.260 1.900 3.540 2.540 ;
        RECT  2.220 1.900 2.500 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.400 0.380 0.820 ;
        RECT  1.140 0.400 1.420 0.820 ;
        RECT  2.180 0.400 2.460 0.820 ;
        RECT  3.180 0.620 3.540 0.820 ;
        RECT  0.100 0.660 3.540 0.820 ;
        RECT  6.340 1.540 8.700 1.740 ;
        RECT  4.260 1.900 4.580 2.100 ;
        RECT  5.260 1.900 5.620 2.100 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  4.260 1.940 6.620 2.100 ;
        RECT  7.380 1.540 7.660 2.100 ;
        RECT  8.420 1.540 8.700 2.100 ;
        RECT  2.660 0.300 8.700 0.460 ;
        RECT  2.660 0.300 3.020 0.500 ;
        RECT  3.700 0.300 4.580 0.500 ;
        RECT  5.260 0.300 5.620 0.500 ;
        RECT  6.300 0.300 6.660 0.500 ;
        RECT  7.340 0.300 7.700 0.500 ;
        RECT  8.380 0.300 8.700 0.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.580 2.400 ;
        RECT  0.000 1.350 1.880 2.400 ;
        RECT  4.110 1.290 8.800 2.400 ;
        RECT  4.130 1.140 8.800 2.400 ;
        RECT  0.000 1.360 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
        RECT  1.580 0.000 4.130 1.290 ;
        RECT  1.580 0.000 4.110 1.350 ;
        RECT  1.880 0.000 4.110 1.360 ;
    END
END OAI211M8HM

MACRO OAI211M4HM
    CLASS CORE ;
    FOREIGN OAI211M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.000 3.500 1.200 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.360 ;
        LAYER ME1 ;
        RECT  3.200 1.000 3.840 1.200 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 1.400 4.300 1.560 ;
        RECT  4.100 1.000 4.300 1.560 ;
        RECT  2.760 0.990 2.920 1.560 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.180 0.900 2.380 1.400 ;
        RECT  0.660 0.900 2.380 1.100 ;
        RECT  0.660 0.900 0.860 1.260 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.240 1.300 1.880 1.500 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.720 4.700 1.880 ;
        RECT  4.500 0.660 4.700 1.880 ;
        RECT  2.860 0.660 4.700 0.820 ;
        RECT  3.900 0.620 4.180 0.820 ;
        RECT  2.860 0.620 3.140 0.820 ;
        RECT  1.980 1.720 2.180 2.030 ;
        RECT  0.860 1.720 1.060 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.260 2.040 4.540 2.540 ;
        RECT  2.500 2.040 2.780 2.540 ;
        RECT  1.380 2.040 1.660 2.540 ;
        RECT  0.340 1.800 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  1.460 -0.140 1.740 0.420 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.400 0.300 4.700 0.460 ;
        RECT  3.380 0.300 3.660 0.500 ;
        RECT  4.420 0.300 4.700 0.500 ;
        RECT  0.640 0.390 0.800 0.740 ;
        RECT  2.400 0.300 2.560 0.740 ;
        RECT  0.640 0.580 2.560 0.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OAI211M4HM

MACRO OAI211M2HM
    CLASS CORE ;
    FOREIGN OAI211M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.890 2.300 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.980 1.540 1.560 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.400 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.480 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.623  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.640 1.720 2.300 1.920 ;
        RECT  1.700 0.620 1.900 1.920 ;
        RECT  1.500 0.620 1.900 0.820 ;
        RECT  0.640 1.560 0.840 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.180 -0.140 0.380 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.980 0.300 2.260 0.460 ;
        RECT  0.980 0.300 1.260 0.540 ;
        RECT  2.060 0.300 2.260 0.600 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END OAI211M2HM

MACRO OAI211M1HM
    CLASS CORE ;
    FOREIGN OAI211M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.890 2.300 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.980 1.540 1.560 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.780 1.100 1.450 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.480 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.540  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.580 1.720 2.300 1.920 ;
        RECT  1.700 0.620 1.900 1.920 ;
        RECT  1.500 0.620 1.900 0.820 ;
        RECT  0.580 1.610 0.860 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.140 0.420 0.500 0.620 ;
        RECT  0.300 -0.140 0.500 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.980 0.300 2.260 0.460 ;
        RECT  0.980 0.300 1.260 0.620 ;
        RECT  2.060 0.300 2.260 0.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END OAI211M1HM

MACRO OAI211M0HM
    CLASS CORE ;
    FOREIGN OAI211M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.890 2.300 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.980 1.540 1.560 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.690 1.100 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.480 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.375  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.580 1.720 2.300 1.920 ;
        RECT  1.700 0.620 1.900 1.920 ;
        RECT  1.500 0.620 1.900 0.820 ;
        RECT  0.580 1.520 0.860 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        RECT  0.100 2.080 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.140 0.420 0.500 0.620 ;
        RECT  0.300 -0.140 0.500 0.620 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END OAI211M0HM

MACRO OAI211B100M8HM
    CLASS CORE ;
    FOREIGN OAI211B100M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.040 4.700 1.240 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  3.720 0.980 5.200 1.300 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.499  LAYER ME1  ;
        ANTENNAGATEAREA 0.499  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.531  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.040 7.100 1.240 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.360 1.020 7.470 1.380 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.580 1.020 9.900 1.640 ;
        RECT  8.200 1.020 9.900 1.280 ;
        END
    END C
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.600 1.240 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.100 1.540 9.380 1.790 ;
        RECT  3.760 1.540 9.380 1.740 ;
        RECT  8.060 1.540 8.340 2.020 ;
        RECT  6.980 1.540 7.260 2.020 ;
        RECT  5.940 1.540 6.220 2.020 ;
        RECT  5.700 0.660 5.900 1.740 ;
        RECT  1.680 0.660 5.900 0.820 ;
        RECT  4.800 0.620 5.160 0.820 ;
        RECT  3.760 0.620 4.120 0.820 ;
        RECT  2.720 0.620 3.080 0.820 ;
        RECT  1.680 0.620 2.040 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.620 1.840 9.900 2.540 ;
        RECT  8.580 1.900 8.860 2.540 ;
        RECT  7.500 1.900 7.780 2.540 ;
        RECT  6.460 1.900 6.740 2.540 ;
        RECT  2.760 1.900 3.040 2.540 ;
        RECT  1.720 1.900 2.000 2.540 ;
        RECT  0.200 1.540 0.480 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.100 -0.140 9.380 0.500 ;
        RECT  8.060 -0.140 8.340 0.500 ;
        RECT  0.200 -0.140 0.480 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.760 0.370 0.960 2.100 ;
        RECT  0.760 1.040 3.120 1.240 ;
        RECT  0.760 1.040 1.000 2.100 ;
        RECT  1.200 1.540 3.520 1.740 ;
        RECT  3.320 1.540 3.520 2.100 ;
        RECT  4.280 1.900 4.640 2.100 ;
        RECT  1.200 1.540 1.480 2.100 ;
        RECT  2.240 1.540 2.520 2.100 ;
        RECT  5.320 1.900 5.640 2.100 ;
        RECT  3.320 1.940 5.640 2.100 ;
        RECT  1.200 0.300 7.300 0.460 ;
        RECT  2.200 0.300 2.560 0.500 ;
        RECT  3.240 0.300 3.600 0.500 ;
        RECT  4.280 0.300 4.640 0.500 ;
        RECT  5.320 0.300 6.260 0.500 ;
        RECT  6.940 0.300 7.300 0.500 ;
        RECT  1.200 0.300 1.480 0.560 ;
        RECT  6.420 0.640 6.770 0.840 ;
        RECT  7.520 0.560 7.800 0.840 ;
        RECT  8.580 0.560 8.860 0.840 ;
        RECT  9.620 0.560 9.900 0.840 ;
        RECT  6.420 0.660 9.900 0.840 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.790 2.400 ;
        RECT  7.930 1.140 10.000 2.400 ;
        RECT  0.000 1.360 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  5.790 0.000 7.930 1.360 ;
    END
END OAI211B100M8HM

MACRO OAI211B100M4HM
    CLASS CORE ;
    FOREIGN OAI211B100M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        ANTENNAGATEAREA 0.244  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.092  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 0.980 4.300 1.180 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.880 0.980 4.560 1.280 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.642  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 0.980 2.300 1.180 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.920 0.980 2.560 1.280 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.460 1.440 5.120 1.600 ;
        RECT  4.900 1.180 5.120 1.600 ;
        RECT  3.460 0.980 3.620 1.600 ;
        END
    END B
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.140 0.500 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.084  LAYER ME1  ;
        ANTENNADIFFAREA 1.084  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.760 3.900 1.960 ;
        LAYER ME2 ;
        RECT  3.700 1.300 3.900 2.020 ;
        LAYER ME1 ;
        RECT  2.040 1.760 4.980 1.920 ;
        RECT  3.500 1.760 3.960 1.960 ;
        RECT  3.140 0.660 3.300 1.920 ;
        RECT  1.540 0.660 3.300 0.820 ;
        RECT  2.580 0.620 2.940 0.820 ;
        RECT  1.540 0.620 1.900 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.220 2.080 5.500 2.540 ;
        RECT  4.100 2.080 4.380 2.540 ;
        RECT  2.980 2.080 3.260 2.540 ;
        RECT  1.260 1.780 1.540 2.540 ;
        RECT  0.100 1.760 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  4.060 -0.140 4.420 0.500 ;
        RECT  0.660 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.700 ;
        RECT  0.100 0.540 0.840 0.700 ;
        RECT  1.480 1.000 1.640 1.600 ;
        RECT  2.820 0.980 2.980 1.600 ;
        RECT  0.680 1.440 2.980 1.600 ;
        RECT  0.680 0.540 0.840 2.100 ;
        RECT  1.180 0.300 3.800 0.460 ;
        RECT  2.060 0.300 2.420 0.500 ;
        RECT  3.100 0.300 3.800 0.500 ;
        RECT  3.640 0.300 3.800 0.820 ;
        RECT  4.980 0.360 5.260 0.820 ;
        RECT  3.640 0.660 5.260 0.820 ;
        RECT  1.180 0.300 1.380 0.840 ;
        RECT  1.060 0.560 1.380 0.840 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END OAI211B100M4HM

MACRO OAI211B100M2HM
    CLASS CORE ;
    FOREIGN OAI211B100M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.060 2.140 1.560 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.080 2.740 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.840 3.500 1.360 ;
        END
    END C
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.030 0.700 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.608  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.010 1.720 3.500 1.920 ;
        RECT  2.900 1.680 3.500 1.920 ;
        RECT  2.900 0.660 3.100 1.920 ;
        RECT  1.740 0.660 3.100 0.840 ;
        RECT  1.740 0.620 2.100 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.660 2.080 2.940 2.540 ;
        RECT  1.320 1.440 1.480 2.540 ;
        RECT  0.300 1.740 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  0.300 -0.140 0.500 0.850 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 0.530 1.020 0.810 ;
        RECT  0.860 1.000 1.480 1.280 ;
        RECT  0.860 0.530 1.020 2.050 ;
        RECT  0.820 1.740 1.020 2.050 ;
        RECT  1.260 0.300 2.620 0.460 ;
        RECT  2.260 0.300 2.620 0.500 ;
        RECT  1.260 0.300 1.540 0.610 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI211B100M2HM

MACRO OAI211B100M1HM
    CLASS CORE ;
    FOREIGN OAI211B100M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.140 2.140 1.500 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.080 2.740 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.840 3.500 1.320 ;
        END
    END C
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 0.580 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.506  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 1.750 3.500 2.100 ;
        RECT  2.100 1.760 3.500 1.920 ;
        RECT  2.900 1.750 3.500 1.920 ;
        RECT  2.900 0.660 3.120 1.920 ;
        RECT  1.700 0.660 3.120 0.840 ;
        RECT  2.100 1.760 2.380 2.100 ;
        RECT  1.700 0.620 2.060 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.660 2.080 2.940 2.540 ;
        RECT  1.220 1.700 1.420 2.540 ;
        RECT  0.180 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  0.180 -0.140 0.460 0.810 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.740 1.040 1.460 1.240 ;
        RECT  0.740 0.530 0.940 2.030 ;
        RECT  1.180 0.300 2.620 0.460 ;
        RECT  2.260 0.300 2.620 0.500 ;
        RECT  1.180 0.300 1.460 0.560 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI211B100M1HM

MACRO OAI211B100M0HM
    CLASS CORE ;
    FOREIGN OAI211B100M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.150 2.060 1.560 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.420 1.080 2.700 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.840 3.500 1.360 ;
        END
    END C
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.090 0.500 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 1.750 3.500 2.100 ;
        RECT  2.020 1.750 3.500 1.920 ;
        RECT  2.020 1.720 3.120 1.920 ;
        RECT  2.900 0.660 3.120 1.920 ;
        RECT  1.620 0.660 3.120 0.840 ;
        RECT  2.020 1.720 2.300 2.100 ;
        RECT  1.620 0.620 1.980 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.620 2.080 2.900 2.540 ;
        RECT  1.140 1.740 1.340 2.540 ;
        RECT  0.100 1.720 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  0.100 -0.140 0.380 0.810 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.040 1.380 1.240 ;
        RECT  0.660 0.530 0.860 2.000 ;
        RECT  1.100 0.300 2.560 0.460 ;
        RECT  2.180 0.300 2.560 0.500 ;
        RECT  1.100 0.300 1.380 0.580 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OAI211B100M0HM

MACRO OA33M8HM
    CLASS CORE ;
    FOREIGN OA33M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.503  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.040 4.300 1.240 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.980 0.980 4.400 1.420 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.887  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.040 5.500 1.240 ;
        LAYER ME2 ;
        RECT  5.300 0.840 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.100 0.980 5.880 1.280 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.887  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.040 2.700 1.240 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.320 0.980 2.960 1.420 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.740 1.440 6.400 1.600 ;
        RECT  6.100 1.000 6.400 1.600 ;
        RECT  4.740 1.000 4.940 1.600 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.440 2.140 1.600 ;
        RECT  1.860 1.000 2.140 1.600 ;
        RECT  0.400 1.000 0.700 1.600 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.460 1.440 8.740 2.100 ;
        RECT  8.500 0.420 8.740 2.100 ;
        RECT  7.420 0.660 8.740 0.840 ;
        RECT  8.460 0.420 8.740 0.840 ;
        RECT  7.420 1.440 8.740 1.640 ;
        RECT  7.420 1.440 7.700 2.100 ;
        RECT  7.420 0.420 7.700 0.840 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.887  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.860 0.980 1.640 1.280 ;
        END
    END B3
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.980 1.440 9.260 2.540 ;
        RECT  7.940 1.900 8.220 2.540 ;
        RECT  6.900 1.440 7.180 2.540 ;
        RECT  5.420 2.080 5.700 2.540 ;
        RECT  1.100 2.080 1.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.980 -0.140 9.260 0.740 ;
        RECT  7.940 -0.140 8.220 0.500 ;
        RECT  6.900 -0.140 7.180 0.500 ;
        RECT  2.660 -0.140 3.020 0.500 ;
        RECT  1.620 -0.140 1.980 0.500 ;
        RECT  0.580 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 1.760 2.300 1.920 ;
        RECT  1.940 1.900 3.300 2.100 ;
        RECT  4.540 1.760 6.620 1.920 ;
        RECT  3.500 1.900 4.820 2.100 ;
        RECT  3.250 0.300 6.700 0.460 ;
        RECT  4.340 0.300 4.620 0.500 ;
        RECT  5.380 0.300 5.660 0.500 ;
        RECT  6.420 0.300 6.700 0.500 ;
        RECT  0.100 0.400 0.380 0.820 ;
        RECT  1.140 0.420 1.420 0.820 ;
        RECT  2.180 0.420 2.460 0.820 ;
        RECT  3.250 0.300 3.470 0.820 ;
        RECT  0.100 0.660 3.470 0.820 ;
        RECT  3.640 0.620 4.100 0.820 ;
        RECT  4.860 0.620 5.140 0.820 ;
        RECT  5.900 0.620 6.180 0.820 ;
        RECT  3.640 0.660 7.160 0.820 ;
        RECT  6.980 0.660 7.160 1.240 ;
        RECT  6.980 1.030 8.340 1.240 ;
        RECT  3.640 0.620 3.800 1.740 ;
        RECT  2.460 1.580 4.340 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
    END
END OA33M8HM

MACRO OA33M4HM
    CLASS CORE ;
    FOREIGN OA33M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 1.000 1.910 1.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.140 1.730 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.040 0.720 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.070 1.000 2.340 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.000 2.740 1.740 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.980 3.280 1.560 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.380 0.660 4.700 1.920 ;
        RECT  3.980 1.700 4.700 1.920 ;
        RECT  3.820 0.660 4.700 0.840 ;
        RECT  3.780 1.900 4.180 2.100 ;
        RECT  3.820 0.390 4.100 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.340 2.080 4.660 2.540 ;
        RECT  3.260 2.080 3.540 2.540 ;
        RECT  0.220 1.720 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.340 -0.140 4.620 0.500 ;
        RECT  3.300 -0.140 3.580 0.560 ;
        RECT  2.260 -0.140 2.540 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.300 2.020 0.460 ;
        RECT  0.580 0.300 0.940 0.500 ;
        RECT  1.740 0.300 2.020 0.820 ;
        RECT  2.780 0.350 3.060 0.820 ;
        RECT  1.740 0.660 3.060 0.820 ;
        RECT  0.100 0.350 0.380 0.820 ;
        RECT  1.100 0.620 1.460 0.820 ;
        RECT  0.100 0.660 1.460 0.820 ;
        RECT  3.600 1.000 4.220 1.280 ;
        RECT  3.600 1.000 3.820 1.740 ;
        RECT  1.300 0.620 1.460 2.060 ;
        RECT  3.440 1.580 3.620 1.920 ;
        RECT  2.930 1.760 3.620 1.920 ;
        RECT  1.300 1.900 3.090 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OA33M4HM

MACRO OA33M2HM
    CLASS CORE ;
    FOREIGN OA33M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 1.000 1.940 1.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.140 1.780 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.220 1.120 0.720 1.570 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.020 2.340 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.040 2.740 1.740 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.980 3.280 1.560 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.900 4.300 2.100 ;
        RECT  4.080 0.300 4.300 2.100 ;
        RECT  3.780 0.300 4.300 0.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.260 2.080 3.540 2.540 ;
        RECT  0.260 1.730 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.300 -0.140 3.580 0.560 ;
        RECT  2.260 -0.140 2.540 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.300 2.020 0.460 ;
        RECT  0.580 0.300 0.940 0.500 ;
        RECT  1.740 0.300 2.020 0.820 ;
        RECT  2.780 0.300 3.060 0.820 ;
        RECT  1.740 0.660 3.060 0.820 ;
        RECT  0.100 0.300 0.380 0.820 ;
        RECT  1.100 0.620 1.460 0.820 ;
        RECT  0.100 0.660 1.460 0.820 ;
        RECT  3.700 0.980 3.920 1.740 ;
        RECT  3.460 1.580 3.920 1.740 ;
        RECT  1.300 0.620 1.460 2.060 ;
        RECT  2.920 1.760 3.620 1.920 ;
        RECT  3.460 1.580 3.620 1.920 ;
        RECT  1.300 1.900 3.080 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OA33M2HM

MACRO OA33M1HM
    CLASS CORE ;
    FOREIGN OA33M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.020 2.340 1.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 1.000 1.940 1.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.140 1.780 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.220 1.140 0.720 1.570 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.040 2.740 1.740 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.980 3.280 1.560 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.900 4.300 2.100 ;
        RECT  4.080 0.330 4.300 2.100 ;
        RECT  3.820 0.330 4.300 0.610 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.260 2.080 3.540 2.540 ;
        RECT  0.260 1.730 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.300 -0.140 3.580 0.560 ;
        RECT  2.260 -0.140 2.540 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.300 2.020 0.460 ;
        RECT  0.580 0.300 0.940 0.500 ;
        RECT  1.740 0.300 2.020 0.820 ;
        RECT  2.780 0.300 3.060 0.820 ;
        RECT  1.740 0.660 3.060 0.820 ;
        RECT  0.100 0.300 0.380 0.820 ;
        RECT  1.100 0.620 1.460 0.820 ;
        RECT  0.100 0.660 1.460 0.820 ;
        RECT  3.700 0.980 3.920 1.740 ;
        RECT  3.460 1.580 3.920 1.740 ;
        RECT  1.300 0.620 1.460 2.060 ;
        RECT  2.920 1.760 3.620 1.920 ;
        RECT  3.460 1.580 3.620 1.920 ;
        RECT  1.300 1.900 3.080 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OA33M1HM

MACRO OA33M0HM
    CLASS CORE ;
    FOREIGN OA33M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 1.000 1.940 1.780 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.140 1.780 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.220 0.980 0.720 1.570 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.020 2.340 1.780 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.040 2.740 1.780 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.980 3.540 1.420 ;
        RECT  2.900 0.980 3.160 1.560 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.900 4.300 2.100 ;
        RECT  4.080 0.300 4.300 2.100 ;
        RECT  3.780 0.300 4.300 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.240 2.080 3.620 2.540 ;
        RECT  0.260 1.730 0.720 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.260 -0.140 3.620 0.820 ;
        RECT  2.220 -0.140 2.580 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.300 2.060 0.460 ;
        RECT  0.580 0.300 0.940 0.500 ;
        RECT  1.680 0.300 2.060 0.820 ;
        RECT  2.740 0.300 3.100 0.820 ;
        RECT  1.680 0.660 3.100 0.820 ;
        RECT  0.100 0.300 0.420 0.820 ;
        RECT  1.100 0.620 1.460 0.820 ;
        RECT  0.100 0.660 1.460 0.820 ;
        RECT  3.700 0.980 3.920 1.740 ;
        RECT  3.360 1.580 3.920 1.740 ;
        RECT  3.360 1.580 3.620 1.920 ;
        RECT  2.920 1.760 3.620 1.920 ;
        RECT  1.300 0.620 1.460 2.100 ;
        RECT  2.920 1.760 3.080 2.100 ;
        RECT  1.300 1.940 3.080 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OA33M0HM

MACRO OA32M8HM
    CLASS CORE ;
    FOREIGN OA32M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.040 2.700 1.240 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.400 0.980 3.040 1.300 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.642  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.040 4.700 1.240 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  4.240 0.980 4.880 1.280 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        ANTENNAGATEAREA 0.278  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.830  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.040 0.980 1.720 1.280 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 1.440 5.400 1.600 ;
        RECT  5.200 1.000 5.400 1.600 ;
        RECT  3.700 0.980 3.960 1.600 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.278  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.440 2.100 1.600 ;
        RECT  1.880 0.980 2.100 1.600 ;
        RECT  0.440 1.000 0.760 1.600 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.700 0.660 7.900 1.650 ;
        RECT  7.500 1.440 7.780 2.100 ;
        RECT  6.460 0.660 7.900 0.860 ;
        RECT  7.500 0.390 7.780 0.860 ;
        RECT  6.460 1.440 7.900 1.640 ;
        RECT  6.460 1.440 6.740 2.100 ;
        RECT  6.460 0.390 6.740 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  8.060 1.480 8.260 2.540 ;
        RECT  6.980 1.900 7.260 2.540 ;
        RECT  5.940 1.440 6.220 2.540 ;
        RECT  4.460 2.080 4.740 2.540 ;
        RECT  1.180 2.080 1.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  8.060 -0.140 8.260 0.720 ;
        RECT  6.980 -0.140 7.260 0.500 ;
        RECT  5.940 -0.140 6.220 0.500 ;
        RECT  1.740 -0.140 2.020 0.500 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.580 1.760 5.660 1.920 ;
        RECT  2.580 1.860 3.860 2.060 ;
        RECT  2.260 0.300 5.740 0.460 ;
        RECT  3.340 0.300 3.620 0.500 ;
        RECT  4.420 0.300 4.700 0.500 ;
        RECT  5.460 0.300 5.740 0.500 ;
        RECT  0.180 0.380 0.460 0.820 ;
        RECT  1.210 0.380 1.500 0.820 ;
        RECT  2.260 0.300 2.540 0.820 ;
        RECT  0.180 0.660 2.540 0.820 ;
        RECT  2.740 0.620 3.100 0.820 ;
        RECT  3.860 0.620 4.220 0.820 ;
        RECT  4.900 0.620 5.260 0.820 ;
        RECT  2.740 0.660 6.170 0.820 ;
        RECT  6.010 0.660 6.170 1.240 ;
        RECT  6.010 1.040 7.480 1.240 ;
        RECT  2.260 1.520 3.420 1.680 ;
        RECT  3.260 0.660 3.420 1.700 ;
        RECT  3.060 1.520 3.420 1.700 ;
        RECT  2.260 1.520 2.420 1.920 ;
        RECT  0.260 1.760 2.420 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END OA32M8HM

MACRO OA32M4HM
    CLASS CORE ;
    FOREIGN OA32M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 1.000 1.900 1.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.000 1.100 1.710 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.090 0.620 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.000 2.300 1.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.110 3.160 1.500 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 1.510 4.700 1.740 ;
        RECT  4.440 0.660 4.700 1.740 ;
        RECT  3.700 0.660 4.700 0.840 ;
        RECT  3.700 1.510 3.980 2.100 ;
        RECT  3.700 0.370 3.980 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.220 1.900 4.500 2.540 ;
        RECT  2.780 1.980 3.420 2.540 ;
        RECT  0.100 1.720 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.220 -0.140 4.500 0.500 ;
        RECT  3.180 -0.140 3.460 0.650 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.300 1.940 0.460 ;
        RECT  0.580 0.300 0.940 0.500 ;
        RECT  1.660 0.300 1.940 0.840 ;
        RECT  2.700 0.370 2.980 0.840 ;
        RECT  1.660 0.680 2.980 0.840 ;
        RECT  0.100 0.370 0.380 0.840 ;
        RECT  1.100 0.620 1.420 0.840 ;
        RECT  0.100 0.680 1.420 0.840 ;
        RECT  3.320 1.020 4.160 1.240 ;
        RECT  3.320 1.020 3.480 1.820 ;
        RECT  2.460 1.660 3.480 1.820 ;
        RECT  1.260 0.620 1.420 2.100 ;
        RECT  2.460 1.660 2.620 2.100 ;
        RECT  1.260 1.870 2.620 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OA32M4HM

MACRO OA32M2HM
    CLASS CORE ;
    FOREIGN OA32M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.960 1.000 3.560 1.500 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.040 2.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.100 1.220 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.680 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.300 1.020 2.760 1.500 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.390 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.060 1.980 3.740 2.540 ;
        RECT  0.180 1.730 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.500 -0.140 3.780 0.710 ;
        RECT  2.500 -0.140 2.780 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.700 0.300 2.220 0.460 ;
        RECT  1.940 0.300 2.220 0.820 ;
        RECT  3.020 0.300 3.290 0.820 ;
        RECT  1.940 0.660 3.290 0.820 ;
        RECT  0.180 0.320 0.460 0.840 ;
        RECT  1.340 0.620 1.620 0.840 ;
        RECT  0.180 0.680 1.620 0.840 ;
        RECT  3.720 0.960 3.920 1.820 ;
        RECT  2.730 1.660 3.920 1.820 ;
        RECT  1.380 0.620 1.540 2.060 ;
        RECT  2.730 1.660 2.890 2.060 ;
        RECT  1.380 1.900 2.890 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OA32M2HM

MACRO OA32M1HM
    CLASS CORE ;
    FOREIGN OA32M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.960 1.000 3.560 1.500 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.000 2.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.000 1.220 1.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.160 0.680 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.300 1.000 2.760 1.500 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.320 4.300 2.090 ;
        RECT  4.020 0.320 4.300 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.060 1.980 3.740 2.540 ;
        RECT  0.180 1.730 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.500 -0.140 3.780 0.600 ;
        RECT  2.500 -0.140 2.780 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.300 2.220 0.460 ;
        RECT  1.940 0.300 2.220 0.840 ;
        RECT  3.020 0.300 3.300 0.840 ;
        RECT  1.940 0.680 3.300 0.840 ;
        RECT  0.180 0.320 0.460 0.840 ;
        RECT  1.260 0.620 1.640 0.840 ;
        RECT  0.180 0.680 1.640 0.840 ;
        RECT  3.720 0.860 3.920 1.820 ;
        RECT  2.730 1.660 3.920 1.820 ;
        RECT  1.380 0.620 1.540 2.060 ;
        RECT  2.730 1.660 2.890 2.060 ;
        RECT  1.380 1.900 2.890 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OA32M1HM

MACRO OA32M0HM
    CLASS CORE ;
    FOREIGN OA32M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.960 1.010 3.560 1.500 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.010 2.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.010 1.220 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.140 0.640 1.560 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.300 1.010 2.760 1.500 ;
        RECT  2.300 1.010 2.570 1.560 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.300 4.300 2.090 ;
        RECT  4.020 0.300 4.300 0.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.060 1.980 3.780 2.540 ;
        RECT  0.180 1.730 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.500 -0.140 3.780 0.600 ;
        RECT  2.500 -0.140 2.780 0.530 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.700 0.300 2.220 0.460 ;
        RECT  1.940 0.300 2.220 0.850 ;
        RECT  2.980 0.300 3.290 0.850 ;
        RECT  1.940 0.690 3.290 0.850 ;
        RECT  0.180 0.320 0.460 0.850 ;
        RECT  0.180 0.620 1.620 0.850 ;
        RECT  3.720 0.930 3.920 1.820 ;
        RECT  2.730 1.660 3.920 1.820 ;
        RECT  1.380 0.620 1.540 2.060 ;
        RECT  2.730 1.660 2.890 2.060 ;
        RECT  1.380 1.900 2.890 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END OA32M0HM

MACRO OA31M8HM
    CLASS CORE ;
    FOREIGN OA31M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER ME1  ;
        ANTENNAGATEAREA 0.274  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.091  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.860 0.980 3.560 1.380 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER ME1  ;
        ANTENNAGATEAREA 0.274  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.167  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.000 1.500 1.200 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.920 0.940 1.740 1.260 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.420 2.240 1.580 ;
        RECT  1.960 0.940 2.240 1.580 ;
        RECT  0.440 0.980 0.760 1.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.790 0.660 7.100 1.380 ;
        RECT  6.700 1.420 6.980 2.100 ;
        RECT  6.790 0.390 6.980 2.100 ;
        RECT  5.660 0.660 7.100 0.860 ;
        RECT  6.700 0.390 6.980 0.860 ;
        RECT  5.660 1.420 6.980 1.640 ;
        RECT  5.660 1.420 5.940 2.100 ;
        RECT  5.660 0.390 5.940 0.860 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.206  LAYER ME1  ;
        ANTENNAGATEAREA 0.206  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.124  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.040 4.300 1.240 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.760 0.980 4.600 1.380 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  7.220 1.540 7.500 2.540 ;
        RECT  6.180 1.900 6.460 2.540 ;
        RECT  5.140 1.480 5.420 2.540 ;
        RECT  4.140 1.860 4.420 2.540 ;
        RECT  1.220 2.060 1.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.220 -0.140 7.500 0.500 ;
        RECT  6.180 -0.140 6.460 0.500 ;
        RECT  5.140 -0.140 5.420 0.710 ;
        RECT  4.140 -0.140 4.420 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 1.740 2.380 1.900 ;
        RECT  0.240 1.740 0.520 2.000 ;
        RECT  2.100 1.900 3.420 2.060 ;
        RECT  0.100 0.300 3.900 0.460 ;
        RECT  0.100 0.300 0.340 0.620 ;
        RECT  3.620 0.300 3.900 0.820 ;
        RECT  4.660 0.300 4.940 0.820 ;
        RECT  3.620 0.660 4.940 0.820 ;
        RECT  0.560 0.620 3.400 0.780 ;
        RECT  4.820 1.020 6.600 1.260 ;
        RECT  2.540 0.620 2.700 1.700 ;
        RECT  2.540 1.540 4.980 1.700 ;
        RECT  3.580 1.540 3.940 2.050 ;
        RECT  4.820 1.020 4.980 2.050 ;
        RECT  4.620 1.540 4.980 2.050 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END OA31M8HM

MACRO OA31M4HM
    CLASS CORE ;
    FOREIGN OA31M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        ANTENNAGATEAREA 0.115  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.559  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.090 2.300 1.290 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.660 1.010 2.300 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 1.010 1.500 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.010 1.100 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.600 1.560 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.780 1.450 3.500 1.740 ;
        RECT  3.260 0.690 3.500 1.740 ;
        RECT  2.780 0.690 3.500 0.850 ;
        RECT  2.660 1.900 3.020 2.100 ;
        RECT  2.780 1.450 3.020 2.100 ;
        RECT  2.780 0.300 3.020 0.850 ;
        RECT  2.700 0.300 3.020 0.530 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.180 -0.140 3.500 0.530 ;
        RECT  2.180 -0.140 2.460 0.530 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  0.100 1.720 0.380 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.580 0.300 1.980 0.460 ;
        RECT  0.580 0.300 0.940 0.530 ;
        RECT  1.620 0.300 1.980 0.530 ;
        RECT  0.100 0.550 0.380 0.850 ;
        RECT  1.100 0.620 1.460 0.850 ;
        RECT  0.100 0.690 2.620 0.850 ;
        RECT  2.460 1.010 3.100 1.290 ;
        RECT  2.460 0.690 2.620 1.740 ;
        RECT  1.660 1.540 2.620 1.740 ;
        RECT  1.660 1.540 1.940 2.050 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OA31M4HM

MACRO OA31M2HM
    CLASS CORE ;
    FOREIGN OA31M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 1.040 1.900 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.200 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.040 0.720 1.560 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.000 2.340 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.410 3.100 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  0.260 1.730 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.280 -0.140 2.590 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 2.080 0.500 ;
        RECT  0.140 0.300 0.420 0.840 ;
        RECT  0.140 0.660 2.720 0.840 ;
        RECT  2.520 0.660 2.720 1.920 ;
        RECT  1.640 1.720 2.720 1.920 ;
        RECT  1.640 1.720 1.920 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.920 2.400 ;
        RECT  1.800 1.140 3.200 2.400 ;
        RECT  0.000 1.180 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
        RECT  0.920 0.000 1.800 1.180 ;
    END
END OA31M2HM

MACRO OA31M1HM
    CLASS CORE ;
    FOREIGN OA31M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.420 1.040 1.900 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.200 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.040 0.720 1.570 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.000 2.360 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.300 3.100 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  0.260 1.730 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.280 -0.140 2.590 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 2.080 0.500 ;
        RECT  0.120 0.300 0.440 0.840 ;
        RECT  0.120 0.660 2.720 0.840 ;
        RECT  2.520 0.660 2.720 1.920 ;
        RECT  1.640 1.720 2.720 1.920 ;
        RECT  1.640 1.720 1.920 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.920 2.400 ;
        RECT  1.800 1.140 3.200 2.400 ;
        RECT  0.000 1.180 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
        RECT  0.920 0.000 1.800 1.180 ;
    END
END OA31M1HM

MACRO OA31M0HM
    CLASS CORE ;
    FOREIGN OA31M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.420 1.040 1.900 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.140 1.560 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.040 0.720 1.570 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.000 2.360 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.300 3.100 2.060 ;
        RECT  2.780 0.300 3.100 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  0.260 1.730 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.280 -0.140 2.590 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 2.080 0.500 ;
        RECT  0.140 0.300 0.420 0.840 ;
        RECT  0.140 0.660 2.720 0.840 ;
        RECT  2.520 0.660 2.720 1.920 ;
        RECT  1.640 1.720 2.720 1.920 ;
        RECT  1.640 1.720 1.920 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.920 2.400 ;
        RECT  1.800 1.140 3.200 2.400 ;
        RECT  0.000 1.180 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
        RECT  0.920 0.000 1.800 1.180 ;
    END
END OA31M0HM

MACRO OA22M8HM
    CLASS CORE ;
    FOREIGN OA22M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.782  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.920 0.980 1.640 1.280 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.642  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.040 0.980 3.680 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.440 4.140 1.600 ;
        RECT  3.940 1.000 4.140 1.600 ;
        RECT  2.500 1.000 2.760 1.600 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.480 1.440 2.100 1.600 ;
        RECT  1.820 1.000 2.100 1.600 ;
        RECT  0.480 0.980 0.760 1.600 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.360 0.840 6.700 1.160 ;
        RECT  6.300 1.440 6.580 2.100 ;
        RECT  6.360 0.370 6.580 2.100 ;
        RECT  6.300 0.370 6.580 0.840 ;
        RECT  5.260 1.440 6.580 1.640 ;
        RECT  5.260 0.660 6.580 0.840 ;
        RECT  5.260 1.440 5.540 2.100 ;
        RECT  5.260 0.370 5.540 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.820 1.540 7.100 2.540 ;
        RECT  5.780 1.900 6.060 2.540 ;
        RECT  4.120 2.080 5.020 2.540 ;
        RECT  4.720 1.660 5.020 2.540 ;
        RECT  2.180 2.080 2.460 2.540 ;
        RECT  0.300 1.840 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.820 -0.140 7.100 0.500 ;
        RECT  5.780 -0.140 6.060 0.500 ;
        RECT  4.740 -0.140 5.020 0.560 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.180 0.300 4.540 0.460 ;
        RECT  3.180 0.300 3.540 0.500 ;
        RECT  4.220 0.300 4.540 0.500 ;
        RECT  0.100 0.360 0.380 0.820 ;
        RECT  1.140 0.360 1.420 0.820 ;
        RECT  2.180 0.300 2.460 0.820 ;
        RECT  0.100 0.660 2.460 0.820 ;
        RECT  2.660 0.620 3.020 0.820 ;
        RECT  3.700 0.620 4.060 0.820 ;
        RECT  2.660 0.660 4.500 0.820 ;
        RECT  4.300 1.000 5.920 1.280 ;
        RECT  4.300 0.660 4.500 1.920 ;
        RECT  1.100 1.760 4.500 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END OA22M8HM

MACRO OA22M4HM
    CLASS CORE ;
    FOREIGN OA22M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        ANTENNAGATEAREA 0.143  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.641  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.040 2.300 1.240 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.980 0.980 2.560 1.400 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.020 1.500 1.660 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.020 1.100 1.660 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.600 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.100 1.470 3.900 1.670 ;
        RECT  3.700 0.660 3.900 1.670 ;
        RECT  3.100 0.660 3.900 0.840 ;
        RECT  3.100 1.470 3.380 2.100 ;
        RECT  3.100 0.300 3.380 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.620 1.890 3.900 2.540 ;
        RECT  2.020 1.880 2.900 2.540 ;
        RECT  0.140 1.790 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.620 -0.140 3.900 0.500 ;
        RECT  2.540 -0.140 2.820 0.380 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.300 2.340 0.460 ;
        RECT  2.180 0.300 2.340 0.820 ;
        RECT  0.100 0.300 0.380 0.820 ;
        RECT  1.140 0.300 1.420 0.820 ;
        RECT  0.100 0.660 1.420 0.820 ;
        RECT  2.180 0.580 2.540 0.820 ;
        RECT  1.660 0.620 1.980 0.820 ;
        RECT  2.720 1.000 3.500 1.280 ;
        RECT  2.720 1.000 2.900 1.720 ;
        RECT  1.660 1.560 2.900 1.720 ;
        RECT  1.660 0.620 1.820 2.020 ;
        RECT  1.020 1.820 1.820 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.440 2.400 ;
        RECT  2.610 1.140 4.000 2.400 ;
        RECT  0.000 1.160 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  1.440 0.000 2.610 1.160 ;
    END
END OA22M4HM

MACRO OA22M2HM
    CLASS CORE ;
    FOREIGN OA22M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.875  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.180 2.300 1.380 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.960 ;
        LAYER ME1 ;
        RECT  2.020 1.020 2.470 1.380 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.240 1.540 1.740 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.240 1.140 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.250 1.240 0.700 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.390 3.500 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.120 1.900 2.980 2.540 ;
        RECT  0.220 1.810 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.740 -0.140 2.940 0.640 ;
        RECT  0.660 -0.140 0.940 0.750 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.220 0.300 2.460 0.460 ;
        RECT  2.260 0.300 2.460 0.840 ;
        RECT  0.170 0.470 0.390 1.070 ;
        RECT  1.220 0.300 1.430 1.070 ;
        RECT  0.170 0.910 1.430 1.070 ;
        RECT  1.700 0.620 1.980 0.820 ;
        RECT  2.940 0.980 3.100 1.740 ;
        RECT  1.700 1.580 3.100 1.740 ;
        RECT  1.700 0.620 1.860 2.060 ;
        RECT  1.060 1.900 1.860 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OA22M2HM

MACRO OA22M1HM
    CLASS CORE ;
    FOREIGN OA22M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.995  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.040 2.300 1.240 ;
        LAYER ME2 ;
        RECT  2.100 0.780 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.020 1.020 2.470 1.400 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.080 1.540 1.740 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.060 1.100 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.260 1.080 0.700 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.340 3.500 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  2.020 1.900 2.300 2.540 ;
        RECT  0.220 1.830 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.700 -0.140 2.900 0.380 ;
        RECT  0.660 -0.140 0.940 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.540 0.460 ;
        RECT  0.140 0.300 0.420 0.840 ;
        RECT  1.180 0.300 1.460 0.840 ;
        RECT  0.140 0.680 1.460 0.840 ;
        RECT  2.340 0.300 2.540 0.860 ;
        RECT  1.700 0.620 2.020 0.820 ;
        RECT  2.940 0.830 3.100 1.740 ;
        RECT  1.700 1.580 3.100 1.740 ;
        RECT  1.700 0.620 1.860 2.060 ;
        RECT  1.060 1.900 1.860 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.550 2.400 ;
        RECT  2.750 1.140 3.600 2.400 ;
        RECT  0.000 1.190 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  1.550 0.000 2.750 1.190 ;
    END
END OA22M1HM

MACRO OA22M0HM
    CLASS CORE ;
    FOREIGN OA22M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.875  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.040 2.300 1.240 ;
        LAYER ME2 ;
        RECT  2.100 0.770 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.020 1.040 2.470 1.400 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.010 1.540 1.740 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.010 1.100 1.740 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 1.010 0.700 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.310 3.500 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  2.020 1.900 2.300 2.540 ;
        RECT  0.220 1.830 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.700 -0.140 2.900 0.380 ;
        RECT  0.660 -0.140 0.940 0.530 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.180 0.300 2.540 0.460 ;
        RECT  0.140 0.370 0.420 0.850 ;
        RECT  1.180 0.300 1.460 0.850 ;
        RECT  0.140 0.690 1.460 0.850 ;
        RECT  2.340 0.300 2.540 0.860 ;
        RECT  1.700 0.650 2.020 0.850 ;
        RECT  2.940 1.190 3.100 1.740 ;
        RECT  1.700 1.580 3.100 1.740 ;
        RECT  1.700 0.650 1.860 2.060 ;
        RECT  1.060 1.900 1.860 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.550 2.400 ;
        RECT  2.750 1.140 3.600 2.400 ;
        RECT  0.000 1.200 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  1.550 0.000 2.750 1.200 ;
    END
END OA22M0HM

MACRO OA222M8HM
    CLASS CORE ;
    FOREIGN OA222M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.780 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.040 1.020 3.680 1.280 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.040 5.900 1.240 ;
        LAYER ME2 ;
        RECT  5.700 0.780 5.900 1.560 ;
        LAYER ME1 ;
        RECT  5.600 1.020 6.240 1.280 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.040 1.500 1.240 ;
        LAYER ME2 ;
        RECT  1.300 0.780 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 1.020 1.600 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 2.020 1.600 ;
        RECT  1.860 0.980 2.020 1.600 ;
        RECT  0.500 1.000 0.700 1.600 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.440 4.140 1.600 ;
        RECT  3.940 1.000 4.140 1.600 ;
        RECT  2.500 1.000 2.740 1.600 ;
        END
    END B2
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.140 1.440 6.700 1.600 ;
        RECT  6.500 1.000 6.700 1.600 ;
        RECT  5.140 1.000 5.340 1.600 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.440 1.440 8.700 2.100 ;
        RECT  8.500 0.370 8.700 2.100 ;
        RECT  7.380 0.660 8.700 0.840 ;
        RECT  8.440 0.370 8.700 0.840 ;
        RECT  7.340 1.440 8.700 1.640 ;
        RECT  7.380 0.370 7.580 0.840 ;
        RECT  7.340 1.440 7.560 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.900 1.900 9.180 2.540 ;
        RECT  7.860 1.900 8.140 2.540 ;
        RECT  6.720 2.080 7.000 2.540 ;
        RECT  4.900 2.080 5.180 2.540 ;
        RECT  4.420 2.080 4.700 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        RECT  0.300 1.900 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.900 -0.140 9.180 0.500 ;
        RECT  7.860 -0.140 8.140 0.500 ;
        RECT  6.860 -0.140 7.060 0.650 ;
        RECT  5.780 -0.140 6.060 0.500 ;
        RECT  4.740 -0.140 5.020 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 4.540 0.460 ;
        RECT  1.140 0.300 1.420 0.500 ;
        RECT  2.180 0.300 2.460 0.500 ;
        RECT  3.220 0.300 3.500 0.500 ;
        RECT  4.260 0.300 4.540 0.500 ;
        RECT  0.140 0.300 0.380 0.660 ;
        RECT  2.630 0.620 2.980 0.820 ;
        RECT  3.740 0.620 4.020 0.820 ;
        RECT  5.300 0.380 5.500 0.820 ;
        RECT  6.340 0.380 6.540 0.820 ;
        RECT  2.630 0.660 6.540 0.820 ;
        RECT  0.620 0.620 0.900 0.820 ;
        RECT  1.660 0.620 1.940 0.820 ;
        RECT  0.620 0.660 2.340 0.820 ;
        RECT  7.000 1.040 8.340 1.240 ;
        RECT  2.180 0.660 2.340 1.920 ;
        RECT  7.000 1.040 7.160 1.920 ;
        RECT  1.100 1.760 7.160 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
    END
END OA222M8HM

MACRO OA222M4HM
    CLASS CORE ;
    FOREIGN OA222M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.075  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.040 1.900 1.240 ;
        LAYER ME2 ;
        RECT  1.700 0.780 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.400 0.980 1.900 1.360 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.565  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.040 2.700 1.240 ;
        LAYER ME2 ;
        RECT  2.500 0.780 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.980 2.700 1.360 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 0.960 1.100 1.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.960 0.360 1.580 ;
        END
    END A2
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.660 3.960 0.860 ;
        RECT  3.660 0.660 3.900 1.320 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.450 1.540 5.100 1.740 ;
        RECT  4.900 0.660 5.100 1.740 ;
        RECT  4.340 0.660 5.100 0.860 ;
        RECT  4.240 1.840 4.650 2.040 ;
        RECT  4.450 1.540 4.650 2.040 ;
        RECT  4.340 0.390 4.540 0.860 ;
        END
    END Z
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.866  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.780 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.000 0.980 3.500 1.300 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.820 1.900 5.100 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.820 -0.140 5.100 0.500 ;
        RECT  3.780 -0.140 4.060 0.500 ;
        RECT  2.740 -0.140 3.020 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.500 0.460 ;
        RECT  2.210 0.300 2.500 0.500 ;
        RECT  1.180 0.300 1.380 0.680 ;
        RECT  0.140 0.300 0.340 0.760 ;
        RECT  3.180 0.340 3.580 0.500 ;
        RECT  1.620 0.620 1.980 0.820 ;
        RECT  3.180 0.340 3.340 0.820 ;
        RECT  1.620 0.660 3.340 0.820 ;
        RECT  0.520 0.620 0.940 0.780 ;
        RECT  4.120 1.040 4.700 1.320 ;
        RECT  4.120 1.040 4.280 1.680 ;
        RECT  1.800 1.520 4.280 1.680 ;
        RECT  0.520 0.620 0.680 1.940 ;
        RECT  1.800 1.520 1.960 1.940 ;
        RECT  0.520 1.780 1.960 1.940 ;
        RECT  2.860 1.520 3.140 2.040 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END OA222M4HM

MACRO OA222M2HM
    CLASS CORE ;
    FOREIGN OA222M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 0.940 1.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.990 0.360 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 1.060 1.900 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.060 2.400 1.560 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.100 1.060 3.500 1.560 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.660 3.900 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.390 4.700 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.840 2.040 4.120 2.540 ;
        RECT  2.220 2.040 2.500 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.900 -0.140 4.180 0.500 ;
        RECT  2.860 -0.140 3.140 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 2.500 0.460 ;
        RECT  2.220 0.300 2.500 0.500 ;
        RECT  1.140 0.300 1.420 0.750 ;
        RECT  0.100 0.300 0.360 0.810 ;
        RECT  3.300 0.340 3.700 0.500 ;
        RECT  1.660 0.620 1.940 0.860 ;
        RECT  3.300 0.340 3.460 0.860 ;
        RECT  1.660 0.660 3.460 0.860 ;
        RECT  0.520 0.620 0.940 0.780 ;
        RECT  0.520 0.620 0.680 2.010 ;
        RECT  1.890 1.720 4.300 1.880 ;
        RECT  4.140 0.980 4.300 1.880 ;
        RECT  0.520 1.850 2.050 2.010 ;
        RECT  2.980 1.720 3.180 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OA222M2HM

MACRO OA222M1HM
    CLASS CORE ;
    FOREIGN OA222M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 0.960 1.100 1.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.970 0.360 1.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.480 1.080 1.900 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.080 2.460 1.560 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.120 1.080 3.500 1.560 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.680 3.900 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.340 4.700 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.840 2.080 4.120 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.900 -0.140 4.180 0.520 ;
        RECT  2.860 -0.140 3.140 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.500 0.460 ;
        RECT  2.220 0.300 2.500 0.520 ;
        RECT  0.140 0.300 0.340 0.810 ;
        RECT  1.180 0.300 1.380 0.810 ;
        RECT  3.300 0.360 3.700 0.520 ;
        RECT  1.660 0.620 1.940 0.880 ;
        RECT  3.300 0.360 3.460 0.880 ;
        RECT  1.660 0.680 3.460 0.880 ;
        RECT  0.520 0.620 0.940 0.780 ;
        RECT  0.520 0.620 0.680 2.010 ;
        RECT  1.890 1.760 4.300 1.920 ;
        RECT  4.140 0.830 4.300 1.920 ;
        RECT  0.520 1.850 2.050 2.010 ;
        RECT  2.980 1.760 3.180 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OA222M1HM

MACRO OA222M0HM
    CLASS CORE ;
    FOREIGN OA222M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.000 1.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.360 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 1.000 1.900 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.060 2.400 1.560 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.120 1.060 3.500 1.560 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.840 3.900 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.310 4.700 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.840 2.080 4.120 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        RECT  0.140 1.830 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.900 -0.140 4.180 0.500 ;
        RECT  2.860 -0.140 3.140 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.550 0.460 ;
        RECT  2.160 0.300 2.550 0.500 ;
        RECT  0.140 0.300 0.340 0.840 ;
        RECT  1.180 0.300 1.380 0.840 ;
        RECT  3.300 0.340 3.700 0.500 ;
        RECT  1.660 0.620 1.940 0.820 ;
        RECT  3.300 0.340 3.460 0.820 ;
        RECT  1.660 0.660 3.460 0.820 ;
        RECT  0.520 0.620 0.940 0.780 ;
        RECT  0.520 0.620 0.680 2.050 ;
        RECT  1.890 1.760 4.300 1.920 ;
        RECT  4.140 0.860 4.300 1.920 ;
        RECT  0.520 1.890 2.050 2.050 ;
        RECT  2.980 1.760 3.180 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OA222M0HM

MACRO OA221M8HM
    CLASS CORE ;
    FOREIGN OA221M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        ANTENNAGATEAREA 0.244  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.049  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.180 1.100 1.380 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.520 1.060 1.160 1.380 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.080 2.300 1.280 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.000 1.020 2.640 1.280 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.080 5.100 1.280 ;
        LAYER ME2 ;
        RECT  4.900 0.840 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.640 1.020 5.280 1.280 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.440 5.800 1.600 ;
        RECT  5.600 1.020 5.800 1.600 ;
        RECT  4.100 1.020 4.340 1.600 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 1.440 3.140 1.600 ;
        RECT  2.900 1.020 3.140 1.600 ;
        RECT  1.560 1.020 1.760 1.600 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.100 0.660 8.300 1.740 ;
        RECT  7.940 1.500 8.140 2.100 ;
        RECT  6.900 0.660 8.300 0.860 ;
        RECT  7.940 0.390 8.140 0.860 ;
        RECT  6.860 1.500 8.300 1.700 ;
        RECT  6.900 0.390 7.100 0.860 ;
        RECT  6.860 1.500 7.080 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.300 2.080 6.580 2.540 ;
        RECT  4.860 2.080 5.140 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 0.400 0.420 0.860 ;
        RECT  1.260 0.400 1.460 0.860 ;
        RECT  2.260 0.620 2.540 0.860 ;
        RECT  3.300 0.620 3.580 0.860 ;
        RECT  0.220 0.660 3.580 0.860 ;
        RECT  1.740 0.300 6.140 0.460 ;
        RECT  1.740 0.300 2.020 0.500 ;
        RECT  2.780 0.300 3.060 0.500 ;
        RECT  4.820 0.300 5.100 0.500 ;
        RECT  5.860 0.300 6.140 0.500 ;
        RECT  3.820 0.300 4.020 0.680 ;
        RECT  4.300 0.620 4.580 0.860 ;
        RECT  5.340 0.620 5.620 0.860 ;
        RECT  4.300 0.660 6.700 0.860 ;
        RECT  6.500 1.060 7.940 1.260 ;
        RECT  0.240 1.580 1.300 1.740 ;
        RECT  1.140 1.580 1.300 1.920 ;
        RECT  6.500 0.660 6.700 1.920 ;
        RECT  1.140 1.760 6.700 1.920 ;
        RECT  0.240 1.580 0.400 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END OA221M8HM

MACRO OA221M4HM
    CLASS CORE ;
    FOREIGN OA221M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.970  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.040 0.700 1.240 ;
        LAYER ME2 ;
        RECT  0.500 0.780 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.250 0.980 0.700 1.380 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.900 1.500 1.560 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.600 1.080 3.100 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.040 2.340 1.600 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.680 3.500 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.000 1.540 4.700 1.740 ;
        RECT  4.500 0.680 4.700 1.740 ;
        RECT  3.940 0.680 4.700 0.880 ;
        RECT  3.900 1.900 4.200 2.100 ;
        RECT  4.000 1.540 4.200 2.100 ;
        RECT  3.940 0.410 4.140 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.420 1.900 4.700 2.540 ;
        RECT  3.340 2.080 3.620 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        RECT  0.300 1.540 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.420 -0.140 4.700 0.520 ;
        RECT  3.380 -0.140 3.660 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.620 0.460 ;
        RECT  2.340 0.300 2.620 0.520 ;
        RECT  0.140 0.300 0.340 0.700 ;
        RECT  1.180 0.300 1.380 0.700 ;
        RECT  2.820 0.360 3.180 0.520 ;
        RECT  1.820 0.620 2.100 0.880 ;
        RECT  2.820 0.360 2.980 0.880 ;
        RECT  1.820 0.680 2.980 0.880 ;
        RECT  0.580 0.620 1.020 0.780 ;
        RECT  3.660 1.040 4.300 1.320 ;
        RECT  0.860 0.620 1.020 1.920 ;
        RECT  3.400 1.600 3.820 1.760 ;
        RECT  3.660 1.040 3.820 1.760 ;
        RECT  0.860 1.760 3.560 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END OA221M4HM

MACRO OA221M2HM
    CLASS CORE ;
    FOREIGN OA221M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        ANTENNAGATEAREA 0.091  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.675  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.130 2.300 1.330 ;
        LAYER ME2 ;
        RECT  2.100 0.780 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.100 1.070 2.600 1.390 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.940 1.500 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 1.240 0.700 1.560 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.030 1.940 1.560 ;
        RECT  1.700 0.620 1.900 1.560 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.710 3.100 1.420 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.440 3.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.060 1.900 3.420 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.340 1.770 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.100 -0.140 3.380 0.510 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.340 0.460 ;
        RECT  1.180 0.300 1.380 0.770 ;
        RECT  2.060 0.300 2.340 0.800 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  0.580 0.620 1.020 0.780 ;
        RECT  3.340 0.900 3.500 1.740 ;
        RECT  2.580 1.580 3.500 1.740 ;
        RECT  0.860 0.620 1.020 1.920 ;
        RECT  0.860 1.760 2.820 1.920 ;
        RECT  2.580 1.580 2.820 2.060 ;
        RECT  2.460 1.760 2.820 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.320 2.400 ;
        RECT  2.950 1.140 4.000 2.400 ;
        RECT  0.000 1.230 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  1.320 0.000 2.950 1.230 ;
    END
END OA221M2HM

MACRO OA221M1HM
    CLASS CORE ;
    FOREIGN OA221M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        ANTENNAGATEAREA 0.091  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.675  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.140 2.300 1.340 ;
        LAYER ME2 ;
        RECT  2.100 0.780 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.100 1.080 2.600 1.400 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 1.060 1.500 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.330 1.080 0.700 1.560 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.140 1.940 1.560 ;
        RECT  1.700 0.680 1.900 1.560 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.840 3.100 1.420 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.380 3.900 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.100 1.900 3.380 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.340 1.830 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.100 -0.140 3.380 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.340 0.460 ;
        RECT  2.060 0.300 2.340 0.800 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  1.180 0.300 1.380 0.830 ;
        RECT  0.580 0.620 1.020 0.780 ;
        RECT  3.340 0.770 3.500 1.740 ;
        RECT  2.480 1.580 3.500 1.740 ;
        RECT  0.860 0.620 1.020 1.920 ;
        RECT  0.860 1.760 2.740 1.920 ;
        RECT  2.480 1.580 2.740 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.320 2.400 ;
        RECT  3.000 1.140 4.000 2.400 ;
        RECT  0.000 1.350 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  1.320 0.000 3.000 1.350 ;
    END
END OA221M1HM

MACRO OA221M0HM
    CLASS CORE ;
    FOREIGN OA221M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.940 1.500 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.960 0.700 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.960 2.600 1.280 ;
        RECT  2.100 0.960 2.300 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.020 1.940 1.560 ;
        RECT  1.700 0.720 1.900 1.560 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.760 0.770 3.160 1.300 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.390 3.900 2.000 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.060 1.840 3.420 2.540 ;
        RECT  1.620 2.040 1.900 2.540 ;
        RECT  0.340 1.720 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.100 -0.140 3.380 0.610 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 2.340 0.460 ;
        RECT  0.140 0.300 0.340 0.770 ;
        RECT  1.180 0.300 1.380 0.770 ;
        RECT  2.060 0.300 2.340 0.800 ;
        RECT  0.580 0.620 1.020 0.780 ;
        RECT  3.340 0.810 3.500 1.680 ;
        RECT  2.580 1.520 3.500 1.680 ;
        RECT  0.860 0.620 1.020 1.880 ;
        RECT  0.860 1.720 2.740 1.880 ;
        RECT  2.580 1.520 2.740 2.060 ;
        RECT  2.540 1.720 2.740 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.320 2.400 ;
        RECT  2.950 1.140 4.000 2.400 ;
        RECT  0.000 1.230 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  1.320 0.000 2.950 1.230 ;
    END
END OA221M0HM

MACRO OA21M8HM
    CLASS CORE ;
    FOREIGN OA21M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.636  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.010 0.980 1.680 1.220 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.960 1.120 2.300 1.340 ;
        RECT  0.500 1.400 2.120 1.560 ;
        RECT  1.960 1.120 2.120 1.560 ;
        RECT  0.500 1.040 0.760 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.460 1.240 5.960 1.560 ;
        RECT  5.480 0.390 5.740 2.080 ;
        RECT  4.420 1.500 5.740 1.700 ;
        RECT  5.460 0.660 5.740 1.700 ;
        RECT  4.460 0.660 5.740 0.860 ;
        RECT  4.460 0.390 4.660 0.860 ;
        RECT  4.420 1.500 4.640 2.080 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        ANTENNAGATEAREA 0.235  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.968  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.170 3.500 1.370 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.200 1.120 3.840 1.370 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.980 1.900 6.260 2.540 ;
        RECT  4.940 1.900 5.220 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        RECT  2.180 2.080 2.460 2.540 ;
        RECT  0.300 1.900 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.980 -0.140 6.260 0.500 ;
        RECT  4.940 -0.140 5.220 0.500 ;
        RECT  3.900 -0.140 4.180 0.500 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 2.620 0.460 ;
        RECT  2.340 0.300 2.620 0.640 ;
        RECT  1.220 0.300 1.500 0.500 ;
        RECT  3.220 0.460 3.700 0.640 ;
        RECT  2.340 0.480 3.700 0.640 ;
        RECT  0.100 0.300 0.380 0.690 ;
        RECT  0.620 0.620 1.040 0.820 ;
        RECT  0.620 0.660 2.060 0.820 ;
        RECT  1.780 0.620 2.060 0.820 ;
        RECT  1.900 0.800 4.260 0.960 ;
        RECT  4.060 1.080 5.240 1.280 ;
        RECT  2.460 1.580 4.260 1.740 ;
        RECT  4.060 0.800 4.260 1.740 ;
        RECT  1.180 1.720 2.660 1.880 ;
        RECT  3.420 1.580 3.620 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END OA21M8HM

MACRO OA21M4HM
    CLASS CORE ;
    FOREIGN OA21M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.580 3.100 1.740 ;
        RECT  2.900 0.660 3.100 1.740 ;
        RECT  2.460 0.660 3.100 0.860 ;
        RECT  2.300 1.900 2.660 2.100 ;
        RECT  2.460 1.580 2.660 2.100 ;
        RECT  2.460 0.300 2.660 0.860 ;
        RECT  2.300 0.300 2.660 0.500 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.414  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.120 1.900 1.320 ;
        LAYER ME2 ;
        RECT  1.700 0.780 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.440 1.060 1.900 1.380 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.650  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 0.780 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.280 1.060 0.700 1.380 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.100 1.560 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 1.900 3.100 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.220 1.540 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.500 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 1.540 0.460 ;
        RECT  1.260 0.300 1.540 0.500 ;
        RECT  0.140 0.300 0.420 0.650 ;
        RECT  0.700 0.620 0.980 0.860 ;
        RECT  0.700 0.660 2.260 0.860 ;
        RECT  2.060 1.020 2.700 1.300 ;
        RECT  2.060 0.660 2.260 1.740 ;
        RECT  1.300 1.580 2.260 1.740 ;
        RECT  1.300 1.580 1.500 2.060 ;
        RECT  1.160 1.860 1.500 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OA21M4HM

MACRO OA21M2HM
    CLASS CORE ;
    FOREIGN OA21M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.155  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.120 1.900 1.320 ;
        LAYER ME2 ;
        RECT  1.700 0.780 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.530 1.060 1.900 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.060 1.220 1.340 ;
        RECT  0.900 1.060 1.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.210 0.740 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.480 0.390 2.700 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.380 1.830 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.260 0.300 1.660 0.460 ;
        RECT  1.380 0.300 1.660 0.500 ;
        RECT  0.260 0.300 0.540 0.560 ;
        RECT  0.820 0.620 1.100 0.900 ;
        RECT  0.820 0.740 2.320 0.900 ;
        RECT  2.120 0.740 2.320 1.740 ;
        RECT  1.320 1.580 2.320 1.740 ;
        RECT  1.320 1.580 1.520 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OA21M2HM

MACRO OA21M1HM
    CLASS CORE ;
    FOREIGN OA21M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.931  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.120 1.900 1.320 ;
        LAYER ME2 ;
        RECT  1.700 0.780 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.560 1.060 1.900 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.020 1.220 1.300 ;
        RECT  0.900 1.020 1.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.200 0.740 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.480 0.320 2.700 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.380 1.790 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.260 0.300 1.660 0.460 ;
        RECT  1.380 0.300 1.660 0.500 ;
        RECT  0.260 0.300 0.540 0.560 ;
        RECT  0.820 0.620 1.100 0.860 ;
        RECT  0.820 0.660 2.320 0.860 ;
        RECT  2.120 0.660 2.320 1.740 ;
        RECT  1.280 1.580 2.320 1.740 ;
        RECT  1.280 1.580 1.480 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OA21M1HM

MACRO OA21M0HM
    CLASS CORE ;
    FOREIGN OA21M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        ANTENNAGATEAREA 0.070  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.931  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 0.780 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.560 1.080 1.900 1.400 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.220 1.320 ;
        RECT  0.900 1.040 1.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.200 0.740 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.480 0.300 2.700 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.380 1.840 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.260 0.300 1.660 0.460 ;
        RECT  1.380 0.300 1.660 0.500 ;
        RECT  0.260 0.300 0.540 0.600 ;
        RECT  0.820 0.620 1.100 0.880 ;
        RECT  0.820 0.680 2.320 0.880 ;
        RECT  2.120 0.680 2.320 1.740 ;
        RECT  1.320 1.580 2.320 1.740 ;
        RECT  1.320 1.580 1.520 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END OA21M0HM

MACRO OA211M8HM
    CLASS CORE ;
    FOREIGN OA211M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME2  ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.900  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.180 1.500 1.380 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.080 1.170 1.720 1.420 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.712  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 0.980 3.500 1.180 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.940 0.980 3.720 1.180 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.340 4.140 1.500 ;
        RECT  3.940 1.040 4.140 1.500 ;
        RECT  2.440 1.040 2.760 1.500 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.850 2.160 1.360 ;
        RECT  0.440 0.850 2.160 1.010 ;
        RECT  0.440 0.850 0.760 1.320 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.660 6.700 1.740 ;
        RECT  6.300 1.450 6.580 2.080 ;
        RECT  6.300 0.520 6.560 0.860 ;
        RECT  5.260 1.450 6.700 1.700 ;
        RECT  5.260 0.660 6.700 0.860 ;
        RECT  5.260 1.450 5.540 2.080 ;
        RECT  5.260 0.520 5.540 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.820 1.900 7.100 2.540 ;
        RECT  5.780 1.900 6.060 2.540 ;
        RECT  4.740 1.900 5.020 2.540 ;
        RECT  4.100 1.980 4.380 2.540 ;
        RECT  2.340 1.980 2.620 2.540 ;
        RECT  1.260 1.900 1.540 2.540 ;
        RECT  0.260 1.750 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.820 -0.140 7.100 0.500 ;
        RECT  5.780 -0.140 6.060 0.500 ;
        RECT  4.740 -0.140 5.020 0.500 ;
        RECT  1.220 -0.140 1.500 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.100 0.300 4.580 0.460 ;
        RECT  3.180 0.300 3.540 0.500 ;
        RECT  4.220 0.300 4.580 0.500 ;
        RECT  2.100 0.300 2.430 0.690 ;
        RECT  0.270 0.530 2.430 0.690 ;
        RECT  2.700 0.620 2.980 0.820 ;
        RECT  3.740 0.620 4.020 0.820 ;
        RECT  2.700 0.660 5.060 0.820 ;
        RECT  4.860 1.080 6.340 1.280 ;
        RECT  4.860 0.660 5.060 1.520 ;
        RECT  4.370 1.320 5.060 1.520 ;
        RECT  0.800 1.580 1.930 1.740 ;
        RECT  4.370 1.320 4.570 1.820 ;
        RECT  1.780 1.660 4.570 1.820 ;
        RECT  1.780 1.660 2.060 1.940 ;
        RECT  0.800 1.580 0.960 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END OA211M8HM

MACRO OA211M4HM
    CLASS CORE ;
    FOREIGN OA211M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.551  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.040 1.100 1.240 ;
        LAYER ME2 ;
        RECT  0.900 0.780 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.890 0.940 1.140 1.420 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.410 1.400 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.760 1.660 1.380 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 0.800 2.300 1.380 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.780 1.540 3.500 1.740 ;
        RECT  3.300 0.660 3.500 1.740 ;
        RECT  2.700 0.660 3.500 0.860 ;
        RECT  2.660 1.900 2.980 2.100 ;
        RECT  2.780 1.540 2.980 2.100 ;
        RECT  2.700 0.390 2.900 0.860 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.180 -0.140 3.460 0.500 ;
        RECT  2.140 -0.140 2.420 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.180 1.900 3.460 2.540 ;
        RECT  2.140 1.900 2.420 2.540 ;
        RECT  1.100 1.900 1.380 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.240 0.300 1.540 0.460 ;
        RECT  1.260 0.300 1.540 0.600 ;
        RECT  0.240 0.300 0.400 0.680 ;
        RECT  0.570 0.620 1.020 0.780 ;
        RECT  2.460 1.060 3.120 1.260 ;
        RECT  0.570 0.620 0.730 1.740 ;
        RECT  2.460 1.060 2.620 1.740 ;
        RECT  0.260 1.580 2.620 1.740 ;
        RECT  0.260 1.580 0.540 2.060 ;
        RECT  1.620 1.580 1.900 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END OA211M4HM

MACRO OA211M2HM
    CLASS CORE ;
    FOREIGN OA211M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 1.900 3.100 2.100 ;
        RECT  2.900 0.430 3.100 2.100 ;
        RECT  2.660 0.430 3.100 0.630 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        ANTENNAGATEAREA 0.091  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.162  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.040 1.100 1.240 ;
        LAYER ME2 ;
        RECT  0.900 0.780 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.890 0.940 1.140 1.420 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.410 1.420 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.660 1.290 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 0.840 2.360 1.400 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.140 -0.140 2.420 0.500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.300 1.900 2.580 2.540 ;
        RECT  1.100 1.900 1.380 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.160 0.300 1.580 0.460 ;
        RECT  1.230 0.300 1.580 0.520 ;
        RECT  0.160 0.300 0.320 0.680 ;
        RECT  0.570 0.620 0.980 0.780 ;
        RECT  0.570 0.620 0.730 1.740 ;
        RECT  2.540 1.000 2.700 1.740 ;
        RECT  0.320 1.580 2.700 1.740 ;
        RECT  0.320 1.580 0.480 2.090 ;
        RECT  1.700 1.580 1.980 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OA211M2HM

MACRO OA211M1HM
    CLASS CORE ;
    FOREIGN OA211M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        ANTENNAGATEAREA 0.091  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.162  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.040 1.100 1.240 ;
        LAYER ME2 ;
        RECT  0.900 0.780 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.890 0.940 1.140 1.420 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.410 1.320 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.660 1.300 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 0.840 2.340 1.320 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 1.900 3.100 2.100 ;
        RECT  2.900 0.360 3.100 2.100 ;
        RECT  2.660 0.360 3.100 0.560 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.140 -0.140 2.420 0.500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.300 1.900 2.580 2.540 ;
        RECT  1.100 1.900 1.380 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 1.580 0.460 ;
        RECT  0.100 0.300 0.380 0.580 ;
        RECT  0.570 0.620 0.980 0.780 ;
        RECT  0.570 0.620 0.730 1.740 ;
        RECT  2.540 0.830 2.700 1.740 ;
        RECT  0.260 1.580 2.700 1.740 ;
        RECT  0.260 1.580 0.540 2.050 ;
        RECT  1.700 1.580 1.980 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OA211M1HM

MACRO OA211M0HM
    CLASS CORE ;
    FOREIGN OA211M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        ANTENNAGATEAREA 0.091  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.162  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.040 1.100 1.240 ;
        LAYER ME2 ;
        RECT  0.900 0.780 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.890 0.940 1.140 1.420 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.410 1.270 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.830 1.660 1.300 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 0.840 2.340 1.320 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 1.900 3.100 2.100 ;
        RECT  2.900 0.320 3.100 2.100 ;
        RECT  2.660 0.320 3.100 0.520 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.140 -0.140 2.420 0.560 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.300 1.900 2.580 2.540 ;
        RECT  1.100 1.900 1.380 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 1.580 0.460 ;
        RECT  0.100 0.300 0.380 0.580 ;
        RECT  0.570 0.620 0.980 0.780 ;
        RECT  0.570 0.620 0.730 1.740 ;
        RECT  2.540 0.830 2.700 1.740 ;
        RECT  0.320 1.580 2.700 1.740 ;
        RECT  0.320 1.580 0.480 2.090 ;
        RECT  1.700 1.580 1.980 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END OA211M0HM

MACRO NR4M8HM
    CLASS CORE ;
    FOREIGN NR4M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        ANTENNAGATEAREA 0.893  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.728  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.180 4.700 1.380 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  1.000 1.260 6.680 1.420 ;
        RECT  6.040 1.120 6.680 1.420 ;
        RECT  4.360 1.120 5.000 1.420 ;
        RECT  2.680 1.120 3.320 1.420 ;
        RECT  1.000 1.120 1.640 1.420 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        ANTENNAGATEAREA 0.893  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.728  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  11.300 1.180 11.500 1.380 ;
        LAYER ME2 ;
        RECT  11.300 0.840 11.500 1.560 ;
        LAYER ME1 ;
        RECT  7.840 1.260 13.520 1.420 ;
        RECT  12.880 1.120 13.520 1.420 ;
        RECT  11.200 1.120 11.840 1.420 ;
        RECT  9.520 1.120 10.160 1.420 ;
        RECT  7.840 1.120 8.480 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.700 0.800 13.940 1.420 ;
        RECT  7.420 0.800 13.940 0.960 ;
        RECT  12.040 0.800 12.680 1.100 ;
        RECT  10.360 0.800 11.000 1.100 ;
        RECT  8.680 0.800 9.320 1.100 ;
        RECT  7.420 0.800 7.580 1.340 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.900 0.800 7.100 1.420 ;
        RECT  0.580 0.800 7.100 0.960 ;
        RECT  5.200 0.800 5.840 1.100 ;
        RECT  3.520 0.800 4.160 1.100 ;
        RECT  1.840 0.800 2.480 1.100 ;
        RECT  0.580 0.800 0.740 1.340 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.688  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.980 1.580 14.300 1.740 ;
        RECT  14.100 0.480 14.300 1.740 ;
        RECT  1.660 0.480 14.300 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.400 2.540 ;
        RECT  6.220 1.900 6.500 2.540 ;
        RECT  4.540 1.900 4.820 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.400 0.140 ;
        RECT  13.100 -0.140 13.380 0.320 ;
        RECT  11.980 -0.140 12.260 0.320 ;
        RECT  11.480 -0.140 11.760 0.320 ;
        RECT  10.360 -0.140 10.640 0.320 ;
        RECT  9.860 -0.140 10.140 0.320 ;
        RECT  8.740 -0.140 9.020 0.320 ;
        RECT  8.260 -0.140 8.540 0.320 ;
        RECT  7.120 -0.140 7.400 0.320 ;
        RECT  5.980 -0.140 6.260 0.320 ;
        RECT  5.500 -0.140 5.780 0.320 ;
        RECT  4.380 -0.140 4.660 0.320 ;
        RECT  3.880 -0.140 4.160 0.320 ;
        RECT  2.760 -0.140 3.040 0.320 ;
        RECT  2.260 -0.140 2.540 0.320 ;
        RECT  1.220 -0.140 1.420 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.300 1.580 7.340 1.740 ;
        RECT  7.060 1.580 7.340 2.060 ;
        RECT  7.060 1.900 14.220 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 14.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.400 1.140 ;
    END
END NR4M8HM

MACRO NR4M6HM
    CLASS CORE ;
    FOREIGN NR4M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.705  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.800 1.260 1.000 1.460 ;
        LAYER ME2 ;
        RECT  0.800 0.840 1.100 1.600 ;
        LAYER ME1 ;
        RECT  0.780 1.050 1.020 1.570 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.240 0.600 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.540 1.540 5.900 1.740 ;
        RECT  5.660 0.410 5.900 1.740 ;
        RECT  4.620 0.680 5.900 0.880 ;
        RECT  4.620 0.410 4.820 0.880 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        ANTENNAGATEAREA 0.098  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.122  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.060 2.570 1.260 ;
        LAYER ME2 ;
        RECT  2.370 0.840 2.700 1.600 ;
        LAYER ME1 ;
        RECT  2.250 0.960 2.570 1.420 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        ANTENNAGATEAREA 0.098  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.963  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.820 1.060 2.020 1.260 ;
        LAYER ME2 ;
        RECT  1.700 0.840 2.020 1.600 ;
        LAYER ME1 ;
        RECT  1.820 0.940 2.090 1.420 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.100 1.900 5.380 2.540 ;
        RECT  4.060 1.480 4.340 2.540 ;
        RECT  3.590 1.900 3.870 2.540 ;
        RECT  2.470 1.900 2.750 2.540 ;
        RECT  0.140 1.840 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.380 0.520 ;
        RECT  4.100 -0.140 4.300 0.600 ;
        RECT  0.100 -0.140 0.380 0.770 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.500 0.620 2.230 0.780 ;
        RECT  1.500 0.620 1.660 2.100 ;
        RECT  2.730 1.060 2.950 1.740 ;
        RECT  1.500 1.580 2.950 1.740 ;
        RECT  1.500 1.580 1.760 2.100 ;
        RECT  1.180 0.300 3.330 0.460 ;
        RECT  0.660 0.600 1.340 0.760 ;
        RECT  3.170 0.300 3.330 1.160 ;
        RECT  3.170 0.960 3.490 1.160 ;
        RECT  1.180 0.300 1.340 2.100 ;
        RECT  1.020 1.840 1.340 2.100 ;
        RECT  3.490 0.400 3.870 0.680 ;
        RECT  3.710 1.080 5.460 1.320 ;
        RECT  3.710 0.400 3.870 1.740 ;
        RECT  3.110 1.580 3.870 1.740 ;
        RECT  3.110 1.580 3.310 2.010 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END NR4M6HM

MACRO NR4M4HM
    CLASS CORE ;
    FOREIGN NR4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.705  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.800 1.260 1.000 1.460 ;
        LAYER ME2 ;
        RECT  0.800 0.900 1.100 1.600 ;
        LAYER ME1 ;
        RECT  0.780 1.050 1.020 1.570 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        ANTENNAGATEAREA 0.098  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.016  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.320 1.080 2.520 1.280 ;
        LAYER ME2 ;
        RECT  2.320 0.840 2.700 1.600 ;
        LAYER ME1 ;
        RECT  2.250 0.940 2.530 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.240 0.600 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.260 1.540 5.100 1.740 ;
        RECT  4.840 0.680 5.100 1.740 ;
        RECT  4.340 0.680 5.100 0.880 ;
        RECT  4.340 0.410 4.540 0.880 ;
        END
    END Z
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        ANTENNAGATEAREA 0.098  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.963  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.820 1.060 2.020 1.260 ;
        LAYER ME2 ;
        RECT  1.700 0.840 2.020 1.600 ;
        LAYER ME1 ;
        RECT  1.820 0.940 2.090 1.420 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.820 1.900 5.100 2.540 ;
        RECT  3.590 1.900 3.870 2.540 ;
        RECT  2.470 1.900 2.750 2.540 ;
        RECT  0.140 1.840 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.820 -0.140 5.100 0.520 ;
        RECT  3.740 -0.140 4.020 0.320 ;
        RECT  0.100 -0.140 0.380 0.770 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.500 0.620 2.230 0.780 ;
        RECT  1.500 0.620 1.660 2.100 ;
        RECT  2.730 1.280 2.950 1.740 ;
        RECT  1.500 1.580 2.950 1.740 ;
        RECT  1.500 1.580 1.760 2.100 ;
        RECT  1.180 0.300 3.270 0.460 ;
        RECT  0.660 0.620 1.340 0.780 ;
        RECT  3.110 0.300 3.270 1.350 ;
        RECT  3.110 1.150 3.490 1.350 ;
        RECT  1.180 0.300 1.340 2.100 ;
        RECT  1.020 1.840 1.340 2.100 ;
        RECT  3.430 0.560 3.870 0.840 ;
        RECT  3.710 1.080 4.550 1.320 ;
        RECT  3.710 0.560 3.870 1.740 ;
        RECT  3.110 1.580 3.870 1.740 ;
        RECT  3.110 1.580 3.310 2.010 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END NR4M4HM

MACRO NR4M2HM
    CLASS CORE ;
    FOREIGN NR4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.031  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.120 1.500 1.320 ;
        LAYER ME2 ;
        RECT  1.300 0.780 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.040 1.120 1.680 1.380 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.031  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.120 3.100 1.320 ;
        LAYER ME2 ;
        RECT  2.900 0.780 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.840 1.120 3.480 1.380 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.800 3.900 1.380 ;
        RECT  2.420 0.800 3.900 0.960 ;
        RECT  2.420 0.800 2.580 1.380 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.940 0.800 2.100 1.380 ;
        RECT  0.500 0.800 2.100 0.960 ;
        RECT  0.500 0.800 0.780 1.380 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.720  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.980 1.540 4.300 1.740 ;
        RECT  4.100 0.480 4.300 1.740 ;
        RECT  1.540 0.480 4.300 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  1.220 1.900 1.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.260 -0.140 3.540 0.320 ;
        RECT  2.140 -0.140 2.420 0.320 ;
        RECT  1.100 -0.140 1.300 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 1.540 2.420 1.740 ;
        RECT  2.220 1.540 2.420 2.060 ;
        RECT  0.380 1.540 0.660 1.950 ;
        RECT  2.220 1.900 4.180 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END NR4M2HM

MACRO NR4M1HM
    CLASS CORE ;
    FOREIGN NR4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        ANTENNAGATEAREA 0.115  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.656  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.090 0.700 1.290 ;
        LAYER ME2 ;
        RECT  0.500 0.780 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.250 1.030 0.700 1.390 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.030 2.300 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.450 1.030 1.900 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.030 1.240 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.527  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.140 1.760 2.700 1.960 ;
        RECT  2.500 0.670 2.700 1.960 ;
        RECT  0.740 0.670 2.700 0.870 ;
        RECT  1.860 0.550 2.060 0.870 ;
        RECT  0.740 0.550 0.940 0.870 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.300 1.590 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.420 -0.140 2.700 0.510 ;
        RECT  0.140 -0.140 0.340 0.730 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END NR4M1HM

MACRO NR4M16HM
    CLASS CORE ;
    FOREIGN NR4M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.786  LAYER ME1  ;
        ANTENNAGATEAREA 1.786  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.984  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.180 4.700 1.380 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  0.760 1.260 13.160 1.420 ;
        RECT  12.520 1.120 13.160 1.420 ;
        RECT  10.840 1.120 11.480 1.420 ;
        RECT  9.160 1.120 9.800 1.420 ;
        RECT  7.480 1.120 8.120 1.420 ;
        RECT  5.800 1.120 6.440 1.420 ;
        RECT  4.120 1.120 4.760 1.420 ;
        RECT  2.440 1.120 3.080 1.420 ;
        RECT  0.760 1.120 1.400 1.420 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.786  LAYER ME1  ;
        ANTENNAGATEAREA 1.786  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.984  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  19.700 1.180 19.900 1.380 ;
        LAYER ME2 ;
        RECT  19.700 0.840 19.900 1.560 ;
        LAYER ME1 ;
        RECT  14.320 1.260 26.720 1.420 ;
        RECT  26.080 1.120 26.720 1.420 ;
        RECT  24.400 1.120 25.040 1.420 ;
        RECT  22.720 1.120 23.360 1.420 ;
        RECT  21.040 1.120 21.680 1.420 ;
        RECT  19.360 1.120 20.000 1.420 ;
        RECT  17.680 1.120 18.320 1.420 ;
        RECT  16.000 1.120 16.640 1.420 ;
        RECT  14.320 1.120 14.960 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.786  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  26.900 0.800 27.140 1.380 ;
        RECT  13.900 0.800 27.140 0.960 ;
        RECT  25.240 0.800 25.880 1.100 ;
        RECT  23.560 0.800 24.200 1.100 ;
        RECT  21.880 0.800 22.520 1.100 ;
        RECT  20.200 0.800 20.840 1.100 ;
        RECT  18.520 0.800 19.160 1.100 ;
        RECT  16.840 0.800 17.480 1.100 ;
        RECT  15.160 0.800 15.800 1.100 ;
        RECT  13.900 0.800 14.060 1.340 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.786  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.420 0.800 13.580 1.340 ;
        RECT  0.100 0.800 13.580 0.960 ;
        RECT  11.680 0.800 12.320 1.100 ;
        RECT  10.000 0.800 10.640 1.100 ;
        RECT  8.320 0.800 8.960 1.100 ;
        RECT  6.640 0.800 7.280 1.100 ;
        RECT  4.960 0.800 5.600 1.100 ;
        RECT  3.280 0.800 3.920 1.100 ;
        RECT  1.600 0.800 2.240 1.100 ;
        RECT  0.100 0.800 0.500 1.380 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.376  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.320 1.580 27.500 1.740 ;
        RECT  27.300 0.480 27.500 1.740 ;
        RECT  1.420 0.480 27.500 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 27.600 2.540 ;
        RECT  12.700 1.900 12.980 2.540 ;
        RECT  11.020 1.900 11.300 2.540 ;
        RECT  9.340 1.900 9.620 2.540 ;
        RECT  7.660 1.900 7.940 2.540 ;
        RECT  5.980 1.900 6.260 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 27.600 0.140 ;
        RECT  26.300 -0.140 26.580 0.320 ;
        RECT  25.180 -0.140 25.460 0.320 ;
        RECT  24.620 -0.140 24.900 0.320 ;
        RECT  23.500 -0.140 23.780 0.320 ;
        RECT  22.940 -0.140 23.220 0.320 ;
        RECT  21.820 -0.140 22.100 0.320 ;
        RECT  21.260 -0.140 21.540 0.320 ;
        RECT  20.140 -0.140 20.420 0.320 ;
        RECT  19.580 -0.140 19.860 0.320 ;
        RECT  18.460 -0.140 18.740 0.320 ;
        RECT  17.960 -0.140 18.240 0.320 ;
        RECT  16.840 -0.140 17.120 0.320 ;
        RECT  16.340 -0.140 16.620 0.320 ;
        RECT  15.220 -0.140 15.500 0.320 ;
        RECT  14.740 -0.140 15.020 0.320 ;
        RECT  13.600 -0.140 13.880 0.320 ;
        RECT  12.460 -0.140 12.740 0.320 ;
        RECT  11.980 -0.140 12.260 0.320 ;
        RECT  10.860 -0.140 11.140 0.320 ;
        RECT  10.360 -0.140 10.640 0.320 ;
        RECT  9.240 -0.140 9.520 0.320 ;
        RECT  8.740 -0.140 9.020 0.320 ;
        RECT  7.620 -0.140 7.900 0.320 ;
        RECT  7.060 -0.140 7.340 0.320 ;
        RECT  5.940 -0.140 6.220 0.320 ;
        RECT  5.380 -0.140 5.660 0.320 ;
        RECT  4.260 -0.140 4.540 0.320 ;
        RECT  3.700 -0.140 3.980 0.320 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.980 -0.140 1.180 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.580 13.930 1.740 ;
        RECT  0.100 1.560 0.440 1.760 ;
        RECT  13.670 1.580 13.930 2.060 ;
        RECT  13.670 1.900 27.500 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 27.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 27.600 1.140 ;
    END
END NR4M16HM

MACRO NR4M12HM
    CLASS CORE ;
    FOREIGN NR4M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.339  LAYER ME1  ;
        ANTENNAGATEAREA 1.339  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.527  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.100 1.140 10.300 1.340 ;
        LAYER ME2 ;
        RECT  10.100 0.780 10.300 1.560 ;
        LAYER ME1 ;
        RECT  10.060 0.800 10.300 1.400 ;
        RECT  0.340 0.800 10.300 0.960 ;
        RECT  8.320 0.800 8.960 1.100 ;
        RECT  6.640 0.800 7.280 1.100 ;
        RECT  4.960 0.800 5.600 1.100 ;
        RECT  3.280 0.800 3.920 1.100 ;
        RECT  1.600 0.800 2.240 1.100 ;
        RECT  0.340 0.800 0.500 1.360 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.339  LAYER ME1  ;
        ANTENNAGATEAREA 1.339  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.759  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  16.100 1.140 16.300 1.340 ;
        LAYER ME2 ;
        RECT  16.100 0.780 16.300 1.560 ;
        LAYER ME1 ;
        RECT  10.960 1.260 19.640 1.420 ;
        RECT  19.360 1.120 19.640 1.420 ;
        RECT  17.680 1.120 18.320 1.420 ;
        RECT  16.000 1.120 16.640 1.420 ;
        RECT  14.320 1.120 14.960 1.420 ;
        RECT  12.640 1.120 13.280 1.420 ;
        RECT  10.960 1.120 11.600 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.339  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  20.100 0.800 20.320 1.400 ;
        RECT  10.540 0.800 20.320 0.960 ;
        RECT  18.520 0.800 19.160 1.100 ;
        RECT  16.840 0.800 17.480 1.100 ;
        RECT  15.160 0.800 15.800 1.100 ;
        RECT  13.480 0.800 14.120 1.100 ;
        RECT  11.800 0.800 12.440 1.100 ;
        RECT  10.540 0.800 10.700 1.360 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.032  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.140 1.580 20.700 1.740 ;
        RECT  20.500 0.480 20.700 1.740 ;
        RECT  1.420 0.480 20.700 0.640 ;
        RECT  19.540 1.580 19.820 1.780 ;
        RECT  17.860 1.580 18.140 1.780 ;
        RECT  16.180 1.580 16.460 1.780 ;
        RECT  14.500 1.580 14.780 1.780 ;
        RECT  12.820 1.580 13.100 1.780 ;
        RECT  11.140 1.580 11.420 1.780 ;
        END
    END Z
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.339  LAYER ME1  ;
        ANTENNAGATEAREA 1.339  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.898  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.170 4.700 1.370 ;
        LAYER ME2 ;
        RECT  4.500 0.780 4.700 1.560 ;
        LAYER ME1 ;
        RECT  0.760 1.260 9.800 1.420 ;
        RECT  9.160 1.120 9.800 1.420 ;
        RECT  7.480 1.120 8.120 1.420 ;
        RECT  5.800 1.120 6.440 1.420 ;
        RECT  4.120 1.120 4.760 1.420 ;
        RECT  2.440 1.120 3.080 1.420 ;
        RECT  0.760 1.120 1.400 1.420 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 20.800 2.540 ;
        RECT  9.340 1.900 9.620 2.540 ;
        RECT  7.660 1.900 7.940 2.540 ;
        RECT  5.980 1.900 6.260 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 20.800 0.140 ;
        RECT  19.580 -0.140 19.860 0.320 ;
        RECT  18.460 -0.140 18.740 0.320 ;
        RECT  17.900 -0.140 18.180 0.320 ;
        RECT  16.780 -0.140 17.060 0.320 ;
        RECT  16.220 -0.140 16.500 0.320 ;
        RECT  15.100 -0.140 15.380 0.320 ;
        RECT  14.600 -0.140 14.880 0.320 ;
        RECT  13.480 -0.140 13.760 0.320 ;
        RECT  12.980 -0.140 13.260 0.320 ;
        RECT  11.860 -0.140 12.140 0.320 ;
        RECT  11.380 -0.140 11.660 0.320 ;
        RECT  10.240 -0.140 10.520 0.320 ;
        RECT  9.100 -0.140 9.380 0.320 ;
        RECT  8.620 -0.140 8.900 0.320 ;
        RECT  7.500 -0.140 7.780 0.320 ;
        RECT  7.000 -0.140 7.280 0.320 ;
        RECT  5.880 -0.140 6.160 0.320 ;
        RECT  5.380 -0.140 5.660 0.320 ;
        RECT  4.260 -0.140 4.540 0.320 ;
        RECT  3.700 -0.140 3.980 0.320 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.980 -0.140 1.180 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.580 10.540 1.740 ;
        RECT  0.100 1.580 0.380 1.900 ;
        RECT  10.340 1.580 10.540 2.100 ;
        RECT  11.980 1.900 12.260 2.100 ;
        RECT  13.660 1.900 13.940 2.100 ;
        RECT  15.340 1.900 15.620 2.100 ;
        RECT  17.020 1.900 17.300 2.100 ;
        RECT  18.700 1.900 18.980 2.100 ;
        RECT  20.380 1.900 20.660 2.100 ;
        RECT  10.340 1.940 20.660 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 20.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 20.800 1.140 ;
    END
END NR4M12HM

MACRO NR4M0HM
    CLASS CORE ;
    FOREIGN NR4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.040 2.300 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 1.040 1.900 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.240 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.040 0.700 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.388  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.900 2.700 2.060 ;
        RECT  2.500 0.680 2.700 2.060 ;
        RECT  0.740 0.680 2.700 0.880 ;
        RECT  1.860 0.540 2.060 0.880 ;
        RECT  0.740 0.540 0.940 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.340 1.800 0.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.420 -0.140 2.700 0.520 ;
        RECT  1.260 -0.140 1.460 0.380 ;
        RECT  0.140 -0.140 0.340 0.820 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END NR4M0HM

MACRO NR4B2M8HM
    CLASS CORE ;
    FOREIGN NR4B2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        ANTENNAGATEAREA 0.893  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.473  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.160 5.100 1.360 ;
        LAYER ME2 ;
        RECT  4.900 1.040 5.100 1.560 ;
        LAYER ME1 ;
        RECT  1.800 1.260 8.380 1.420 ;
        RECT  8.220 0.960 8.380 1.420 ;
        RECT  6.480 1.120 7.120 1.420 ;
        RECT  4.800 1.120 5.440 1.420 ;
        RECT  3.120 1.120 3.760 1.420 ;
        RECT  1.800 1.040 2.080 1.420 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.300 1.120 15.500 1.560 ;
        RECT  8.900 1.260 15.500 1.420 ;
        RECT  15.200 1.120 15.500 1.420 ;
        RECT  13.520 1.120 14.160 1.420 ;
        RECT  11.840 1.120 12.480 1.420 ;
        RECT  10.160 1.120 10.800 1.420 ;
        RECT  8.900 0.900 9.060 1.420 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.900 1.080 1.220 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.900 1.020 17.100 1.560 ;
        RECT  16.200 1.020 17.100 1.340 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.848  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.540 1.580 14.880 1.740 ;
        RECT  2.940 0.480 14.060 0.640 ;
        RECT  8.440 0.480 8.760 0.700 ;
        RECT  8.540 0.480 8.740 1.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.600 2.540 ;
        RECT  16.900 1.900 17.180 2.540 ;
        RECT  15.860 1.900 16.140 2.540 ;
        RECT  7.500 1.900 7.780 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.140 1.900 4.420 2.540 ;
        RECT  2.460 1.900 2.740 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.530 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.600 0.140 ;
        RECT  16.900 -0.140 17.180 0.560 ;
        RECT  15.860 -0.140 16.140 0.500 ;
        RECT  14.580 -0.140 14.860 0.320 ;
        RECT  12.960 -0.140 13.240 0.320 ;
        RECT  11.340 -0.140 12.120 0.320 ;
        RECT  10.220 -0.140 10.500 0.320 ;
        RECT  8.400 -0.140 8.680 0.320 ;
        RECT  6.780 -0.140 7.540 0.320 ;
        RECT  5.160 -0.140 5.940 0.320 ;
        RECT  3.540 -0.140 4.320 0.320 ;
        RECT  2.420 -0.140 2.700 0.320 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        RECT  0.140 -0.140 0.340 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.390 0.860 0.740 ;
        RECT  0.660 0.540 1.460 0.740 ;
        RECT  1.260 0.640 2.480 0.840 ;
        RECT  2.280 0.800 7.960 0.960 ;
        RECT  2.280 0.800 2.920 1.100 ;
        RECT  3.960 0.800 4.600 1.100 ;
        RECT  5.640 0.800 6.280 1.100 ;
        RECT  7.320 0.800 7.960 1.100 ;
        RECT  1.260 0.540 1.460 1.740 ;
        RECT  0.620 1.500 1.460 1.740 ;
        RECT  1.620 1.580 8.160 1.740 ;
        RECT  1.620 1.580 1.900 1.800 ;
        RECT  7.960 1.580 8.160 2.100 ;
        RECT  8.340 1.900 8.620 2.100 ;
        RECT  10.340 1.900 10.620 2.100 ;
        RECT  12.020 1.900 12.300 2.100 ;
        RECT  13.700 1.900 13.980 2.100 ;
        RECT  15.380 1.900 15.660 2.100 ;
        RECT  7.960 1.940 15.660 2.100 ;
        RECT  15.700 0.660 16.660 0.820 ;
        RECT  16.380 0.420 16.660 0.820 ;
        RECT  9.320 0.800 15.900 0.960 ;
        RECT  9.320 0.800 9.960 1.100 ;
        RECT  11.000 0.800 11.640 1.100 ;
        RECT  12.860 0.800 13.140 1.100 ;
        RECT  14.360 0.800 14.640 1.100 ;
        RECT  15.700 0.660 15.900 1.740 ;
        RECT  15.700 1.540 16.620 1.740 ;
        RECT  16.420 1.540 16.620 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 17.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.600 1.140 ;
    END
END NR4B2M8HM

MACRO NR4B2M4HM
    CLASS CORE ;
    FOREIGN NR4B2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.461  LAYER ME1  ;
        ANTENNAGATEAREA 0.461  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.491  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.140 3.100 1.340 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  1.280 1.260 4.500 1.420 ;
        RECT  4.340 1.000 4.500 1.420 ;
        RECT  2.600 1.120 3.240 1.420 ;
        RECT  1.280 1.060 1.560 1.420 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.461  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.100 1.060 8.300 1.560 ;
        RECT  5.020 1.260 8.300 1.420 ;
        RECT  7.960 1.060 8.300 1.420 ;
        RECT  6.280 1.120 6.920 1.420 ;
        RECT  5.020 1.020 5.180 1.420 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 0.840 0.700 1.220 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.900 0.840 9.300 1.220 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.392  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.660 1.580 7.620 1.740 ;
        RECT  2.420 0.480 7.100 0.640 ;
        RECT  4.660 0.480 4.860 1.740 ;
        RECT  4.440 0.480 4.860 0.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.140 1.900 9.420 2.540 ;
        RECT  3.620 1.900 3.900 2.540 ;
        RECT  1.940 1.900 2.220 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.140 -0.140 9.420 0.500 ;
        RECT  7.340 -0.140 7.620 0.500 ;
        RECT  5.740 -0.140 6.500 0.320 ;
        RECT  4.620 -0.140 4.900 0.320 ;
        RECT  3.020 -0.140 3.780 0.320 ;
        RECT  1.940 -0.140 2.220 0.500 ;
        RECT  0.160 -0.140 0.320 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.480 1.100 0.640 ;
        RECT  0.900 0.680 1.960 0.880 ;
        RECT  1.760 0.800 4.080 0.960 ;
        RECT  1.760 0.800 2.400 1.100 ;
        RECT  3.440 0.800 4.080 1.100 ;
        RECT  0.900 0.480 1.100 1.740 ;
        RECT  0.620 1.580 0.900 2.060 ;
        RECT  1.580 1.580 4.300 1.740 ;
        RECT  4.100 1.580 4.300 2.060 ;
        RECT  1.580 1.580 1.740 2.060 ;
        RECT  1.060 1.900 1.740 2.060 ;
        RECT  2.780 1.580 3.060 2.060 ;
        RECT  4.100 1.900 8.460 2.060 ;
        RECT  8.500 0.340 8.940 0.500 ;
        RECT  7.600 0.680 8.700 0.880 ;
        RECT  5.440 0.800 7.760 0.960 ;
        RECT  5.440 0.800 6.080 1.100 ;
        RECT  7.120 0.800 7.760 1.100 ;
        RECT  8.500 0.340 8.700 1.740 ;
        RECT  8.620 1.580 8.900 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
    END
END NR4B2M4HM

MACRO NR4B2M2HM
    CLASS CORE ;
    FOREIGN NR4B2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.840 0.800 5.120 1.100 ;
        RECT  4.900 0.440 5.120 1.100 ;
        RECT  3.720 0.800 5.120 0.960 ;
        RECT  3.580 1.060 3.880 1.340 ;
        RECT  3.720 0.800 3.880 1.340 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.800 3.060 1.340 ;
        RECT  1.520 0.800 3.060 0.960 ;
        RECT  1.700 0.440 1.900 0.960 ;
        RECT  1.520 0.800 1.800 1.100 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 1.040 0.740 1.560 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.840 1.040 6.300 1.320 ;
        RECT  5.900 0.840 6.300 1.320 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.720  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 1.580 4.500 1.740 ;
        RECT  2.580 0.480 4.060 0.640 ;
        RECT  3.220 0.480 3.560 0.700 ;
        RECT  3.220 0.480 3.420 1.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  6.020 1.580 6.300 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  0.340 1.850 0.620 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  6.060 -0.140 6.260 0.640 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.180 -0.140 3.460 0.320 ;
        RECT  2.100 -0.140 2.380 0.500 ;
        RECT  0.360 -0.140 0.580 0.800 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.000 1.120 2.640 1.420 ;
        RECT  0.900 1.260 2.640 1.420 ;
        RECT  0.900 0.520 1.100 2.060 ;
        RECT  1.300 1.580 2.820 1.740 ;
        RECT  2.660 1.580 2.820 2.060 ;
        RECT  2.660 1.900 5.340 2.060 ;
        RECT  5.540 0.360 5.740 0.880 ;
        RECT  5.300 0.680 5.740 0.880 ;
        RECT  4.200 1.120 4.640 1.340 ;
        RECT  4.440 1.260 5.500 1.420 ;
        RECT  5.300 0.680 5.500 1.740 ;
        RECT  5.300 1.580 5.820 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END NR4B2M2HM

MACRO NR4B2M1HM
    CLASS CORE ;
    FOREIGN NR4B2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 1.040 2.300 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.700 1.560 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.900 0.760 1.320 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 1.040 3.900 1.560 ;
        RECT  3.320 1.040 3.900 1.320 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.478  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.900 2.940 2.060 ;
        RECT  2.500 0.680 2.700 2.060 ;
        RECT  2.380 0.560 2.580 0.880 ;
        RECT  1.240 0.680 2.700 0.880 ;
        RECT  1.240 0.560 1.460 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.620 2.080 3.900 2.540 ;
        RECT  0.800 1.900 1.090 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.940 -0.140 3.220 0.520 ;
        RECT  1.740 -0.140 2.020 0.520 ;
        RECT  0.620 -0.140 0.900 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.080 0.740 ;
        RECT  0.920 0.520 1.080 1.700 ;
        RECT  0.920 1.040 1.120 1.700 ;
        RECT  0.160 1.540 1.120 1.700 ;
        RECT  3.580 0.560 3.780 0.880 ;
        RECT  2.860 0.680 3.780 0.880 ;
        RECT  2.860 0.680 3.080 1.740 ;
        RECT  2.860 1.580 3.420 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END NR4B2M1HM

MACRO NR4B2M0HM
    CLASS CORE ;
    FOREIGN NR4B2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 1.040 2.300 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.700 1.560 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.480 0.840 0.760 1.320 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 1.040 3.900 1.560 ;
        RECT  3.320 1.040 3.900 1.320 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.370  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.600 2.840 1.960 ;
        RECT  2.500 0.680 2.700 1.960 ;
        RECT  2.400 0.520 2.560 0.880 ;
        RECT  1.280 0.680 2.700 0.880 ;
        RECT  1.280 0.520 1.440 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.620 1.990 3.900 2.540 ;
        RECT  0.800 1.660 1.090 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.940 -0.140 3.220 0.520 ;
        RECT  1.740 -0.140 2.020 0.320 ;
        RECT  0.620 -0.140 0.900 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.080 0.680 ;
        RECT  0.920 0.520 1.080 1.320 ;
        RECT  0.920 1.040 1.120 1.320 ;
        RECT  0.100 0.520 0.320 1.760 ;
        RECT  0.100 1.540 0.480 1.760 ;
        RECT  3.580 0.560 3.780 0.880 ;
        RECT  2.860 0.680 3.780 0.880 ;
        RECT  2.860 0.680 3.160 1.320 ;
        RECT  3.000 0.680 3.160 1.660 ;
        RECT  3.000 1.500 3.420 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END NR4B2M0HM

MACRO NR4B1M8HM
    CLASS CORE ;
    FOREIGN NR4B1M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        ANTENNAGATEAREA 0.893  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.518  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  10.900 1.160 11.100 1.360 ;
        LAYER ME2 ;
        RECT  10.900 1.040 11.100 1.560 ;
        LAYER ME1 ;
        RECT  9.120 1.260 14.440 1.420 ;
        RECT  14.160 1.120 14.440 1.420 ;
        RECT  12.660 1.120 12.940 1.420 ;
        RECT  10.800 1.120 11.440 1.420 ;
        RECT  9.120 1.120 9.760 1.420 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        ANTENNAGATEAREA 0.893  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.531  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.160 5.100 1.360 ;
        LAYER ME2 ;
        RECT  4.900 1.040 5.100 1.560 ;
        LAYER ME1 ;
        RECT  1.700 1.260 8.380 1.420 ;
        RECT  8.220 0.960 8.380 1.420 ;
        RECT  6.480 1.120 7.120 1.420 ;
        RECT  4.800 1.120 5.440 1.420 ;
        RECT  3.120 1.120 3.760 1.420 ;
        RECT  1.700 1.040 2.020 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.900 0.800 15.120 1.360 ;
        RECT  8.700 0.800 15.120 0.960 ;
        RECT  13.320 0.800 13.960 1.100 ;
        RECT  11.640 0.800 12.280 1.100 ;
        RECT  9.960 0.800 10.600 1.100 ;
        RECT  8.700 0.800 8.860 1.320 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.900 1.080 1.220 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.848  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.300 0.480 15.500 1.740 ;
        RECT  13.140 1.580 15.500 1.740 ;
        RECT  2.940 0.480 15.500 0.640 ;
        RECT  12.300 1.600 13.300 1.760 ;
        RECT  9.260 1.580 12.460 1.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  7.500 1.900 7.780 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.140 1.900 4.420 2.540 ;
        RECT  2.460 1.900 2.740 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.560 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  14.380 -0.140 14.660 0.320 ;
        RECT  12.760 -0.140 13.040 0.320 ;
        RECT  11.140 -0.140 11.920 0.320 ;
        RECT  10.020 -0.140 10.300 0.320 ;
        RECT  8.400 -0.140 8.680 0.320 ;
        RECT  6.780 -0.140 7.540 0.320 ;
        RECT  5.160 -0.140 5.940 0.320 ;
        RECT  3.540 -0.140 4.320 0.320 ;
        RECT  2.420 -0.140 2.700 0.320 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        RECT  0.140 -0.140 0.340 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.390 0.860 0.740 ;
        RECT  0.660 0.540 1.460 0.740 ;
        RECT  1.260 0.640 2.480 0.840 ;
        RECT  2.280 0.800 7.960 0.960 ;
        RECT  2.280 0.800 2.920 1.100 ;
        RECT  3.960 0.800 4.600 1.100 ;
        RECT  5.640 0.800 6.280 1.100 ;
        RECT  7.320 0.800 7.960 1.100 ;
        RECT  1.260 0.540 1.460 1.740 ;
        RECT  0.620 1.500 1.460 1.740 ;
        RECT  1.620 1.580 8.700 1.740 ;
        RECT  1.620 1.580 1.900 1.800 ;
        RECT  8.500 1.580 8.700 2.100 ;
        RECT  10.140 1.900 10.420 2.100 ;
        RECT  11.820 1.900 12.100 2.100 ;
        RECT  13.500 1.900 13.780 2.100 ;
        RECT  15.180 1.900 15.460 2.100 ;
        RECT  8.500 1.940 15.460 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.140 ;
    END
END NR4B1M8HM

MACRO NR4B1M4HM
    CLASS CORE ;
    FOREIGN NR4B1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.796  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.170 5.500 1.370 ;
        LAYER ME2 ;
        RECT  5.300 1.040 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.240 1.260 7.200 1.420 ;
        RECT  6.900 1.120 7.200 1.420 ;
        RECT  5.240 1.120 5.880 1.420 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.694  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.140 1.500 1.340 ;
        LAYER ME2 ;
        RECT  1.300 1.040 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.280 1.260 4.500 1.420 ;
        RECT  4.340 1.000 4.500 1.420 ;
        RECT  2.600 1.120 3.240 1.420 ;
        RECT  1.280 1.010 1.560 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.700 0.800 7.920 1.160 ;
        RECT  4.820 0.800 7.920 0.960 ;
        RECT  6.080 0.800 6.720 1.100 ;
        RECT  4.820 0.800 4.980 1.360 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 0.840 0.700 1.300 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.344  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.380 1.580 8.300 1.740 ;
        RECT  8.100 0.440 8.300 1.740 ;
        RECT  2.420 0.480 8.300 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  3.620 1.900 3.900 2.540 ;
        RECT  1.940 1.900 2.220 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.140 -0.140 7.420 0.320 ;
        RECT  5.660 -0.140 6.300 0.320 ;
        RECT  4.520 -0.140 4.800 0.320 ;
        RECT  3.020 -0.140 3.660 0.320 ;
        RECT  1.940 -0.140 2.220 0.520 ;
        RECT  0.100 -0.140 0.380 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.490 1.100 0.650 ;
        RECT  0.900 0.680 1.920 0.840 ;
        RECT  1.760 0.800 4.080 0.960 ;
        RECT  1.760 0.800 2.400 1.100 ;
        RECT  3.440 0.800 4.080 1.100 ;
        RECT  0.900 0.490 1.100 1.740 ;
        RECT  0.620 1.580 0.900 2.060 ;
        RECT  1.580 1.580 4.260 1.740 ;
        RECT  4.100 1.580 4.260 2.060 ;
        RECT  1.580 1.580 1.740 2.060 ;
        RECT  1.060 1.900 1.740 2.060 ;
        RECT  2.780 1.580 3.060 2.060 ;
        RECT  4.100 1.900 8.260 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END NR4B1M4HM

MACRO NR4B1M2HM
    CLASS CORE ;
    FOREIGN NR4B1M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.009  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.140 3.900 1.340 ;
        LAYER ME2 ;
        RECT  3.700 1.040 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.560 1.120 4.200 1.370 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 0.800 2.820 1.360 ;
        RECT  1.280 0.800 2.820 0.960 ;
        RECT  1.280 0.440 1.560 0.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.460 0.800 4.700 1.400 ;
        RECT  3.140 0.800 4.700 0.960 ;
        RECT  3.140 0.800 3.300 1.360 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.180 0.500 1.560 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.720  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 1.580 5.100 1.740 ;
        RECT  4.900 0.480 5.100 1.740 ;
        RECT  2.260 0.480 5.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  1.940 1.900 2.220 2.540 ;
        RECT  0.100 1.780 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  3.980 -0.140 4.260 0.320 ;
        RECT  2.860 -0.140 3.140 0.320 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        RECT  0.100 -0.140 0.380 0.800 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.760 1.120 2.400 1.420 ;
        RECT  0.660 1.260 2.400 1.420 ;
        RECT  0.660 0.520 0.860 1.980 ;
        RECT  1.060 1.580 2.580 1.740 ;
        RECT  2.420 1.580 2.580 2.060 ;
        RECT  2.420 1.900 4.900 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END NR4B1M2HM

MACRO NR4B1M1HM
    CLASS CORE ;
    FOREIGN NR4B1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.700 1.320 ;
        RECT  1.300 1.040 1.500 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.040 2.300 1.560 ;
        RECT  2.020 1.040 2.300 1.320 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.040 3.100 1.560 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.900 0.760 1.320 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.478  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.900 2.940 2.060 ;
        RECT  2.500 0.680 2.700 2.060 ;
        RECT  2.380 0.560 2.580 0.880 ;
        RECT  1.240 0.680 2.700 0.880 ;
        RECT  1.240 0.560 1.460 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  0.800 1.900 1.090 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.940 -0.140 3.220 0.780 ;
        RECT  1.740 -0.140 2.020 0.320 ;
        RECT  0.620 -0.140 0.900 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.080 0.740 ;
        RECT  0.920 0.520 1.080 1.700 ;
        RECT  0.920 1.040 1.120 1.700 ;
        RECT  0.160 1.540 1.120 1.700 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END NR4B1M1HM

MACRO NR4B1M0HM
    CLASS CORE ;
    FOREIGN NR4B1M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.700 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.020 1.040 2.300 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.040 2.720 1.560 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.480 0.840 0.760 1.320 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.396  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.720 3.100 1.960 ;
        RECT  2.900 0.680 3.100 1.960 ;
        RECT  1.280 0.680 3.100 0.840 ;
        RECT  2.300 0.560 2.580 0.840 ;
        RECT  1.280 0.560 1.500 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  0.800 1.660 1.090 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.340 ;
        RECT  1.700 -0.140 1.980 0.320 ;
        RECT  0.620 -0.140 0.900 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.520 1.080 0.680 ;
        RECT  0.920 0.520 1.080 1.320 ;
        RECT  0.920 1.040 1.120 1.320 ;
        RECT  0.100 0.520 0.320 1.760 ;
        RECT  0.100 1.540 0.480 1.760 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END NR4B1M0HM

MACRO NR3M8HM
    CLASS CORE ;
    FOREIGN NR3M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.476  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.300 1.080 5.900 1.280 ;
        RECT  5.700 0.840 5.900 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.476  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.800 3.500 1.340 ;
        RECT  0.340 0.800 3.500 0.960 ;
        RECT  1.600 0.800 2.240 1.040 ;
        RECT  0.340 0.800 0.500 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.476  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.240 3.080 1.400 ;
        RECT  2.440 1.120 3.080 1.400 ;
        RECT  1.700 1.240 1.900 1.560 ;
        RECT  0.760 1.120 1.160 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.294  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 1.580 5.340 1.740 ;
        RECT  3.900 0.680 5.300 0.880 ;
        RECT  5.020 0.340 5.300 0.880 ;
        RECT  3.980 0.340 4.300 0.880 ;
        RECT  3.900 0.480 4.100 1.740 ;
        RECT  0.620 0.480 4.300 0.640 ;
        RECT  2.860 0.420 3.140 0.640 ;
        RECT  1.740 0.420 2.020 0.640 ;
        RECT  0.620 0.420 0.900 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.540 -0.140 5.820 0.500 ;
        RECT  4.500 -0.140 4.780 0.500 ;
        RECT  3.420 -0.140 3.700 0.320 ;
        RECT  2.300 -0.140 2.580 0.320 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        RECT  0.140 -0.140 0.340 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.580 1.540 1.740 ;
        RECT  2.300 1.580 3.260 1.740 ;
        RECT  0.100 1.580 0.380 1.840 ;
        RECT  1.380 1.580 1.540 2.060 ;
        RECT  3.100 1.580 3.260 2.060 ;
        RECT  2.300 1.580 2.460 2.060 ;
        RECT  1.380 1.900 2.460 2.060 ;
        RECT  3.100 1.900 5.860 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END NR3M8HM

MACRO NR3M6HM
    CLASS CORE ;
    FOREIGN NR3M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.358  LAYER ME1  ;
        ANTENNAGATEAREA 0.358  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.036  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.140 2.700 1.340 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.080 1.080 3.160 1.400 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.358  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.640 1.080 4.720 1.320 ;
        RECT  4.500 0.840 4.720 1.320 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.358  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.080 1.600 1.400 ;
        RECT  0.500 1.080 0.700 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.111  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.580 5.100 2.060 ;
        RECT  4.900 0.340 5.100 2.060 ;
        RECT  4.820 0.340 5.100 0.560 ;
        RECT  3.320 1.580 5.100 1.740 ;
        RECT  0.660 0.680 4.060 0.880 ;
        RECT  3.780 0.340 4.060 0.880 ;
        RECT  3.320 0.680 3.480 1.740 ;
        RECT  2.740 0.340 3.020 0.880 ;
        RECT  1.700 0.340 1.980 0.880 ;
        RECT  0.660 0.340 0.940 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.140 1.900 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.300 -0.140 4.580 0.500 ;
        RECT  3.260 -0.140 3.540 0.500 ;
        RECT  2.220 -0.140 2.500 0.500 ;
        RECT  1.180 -0.140 1.460 0.500 ;
        RECT  0.180 -0.140 0.380 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.860 1.580 3.060 1.740 ;
        RECT  0.860 1.580 1.020 2.060 ;
        RECT  0.620 1.900 1.020 2.060 ;
        RECT  1.700 1.580 1.980 2.060 ;
        RECT  2.180 1.900 4.620 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END NR3M6HM

MACRO NR3M4HM
    CLASS CORE ;
    FOREIGN NR3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.918  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.580 1.140 1.780 1.340 ;
        LAYER ME2 ;
        RECT  1.580 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.280 1.120 1.880 1.370 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.080 1.120 2.400 1.320 ;
        RECT  0.760 1.580 2.280 1.740 ;
        RECT  2.080 1.120 2.280 1.740 ;
        RECT  0.760 1.120 1.100 1.740 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.620 0.800 2.780 1.260 ;
        RECT  0.100 0.800 2.780 0.960 ;
        RECT  0.100 0.800 0.500 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.686  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.520 3.100 1.680 ;
        RECT  2.940 0.420 3.100 1.680 ;
        RECT  1.660 0.480 3.100 0.640 ;
        RECT  2.820 0.420 3.100 0.640 ;
        RECT  1.380 1.900 2.700 2.060 ;
        RECT  2.500 1.520 2.700 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.880 1.840 3.100 2.540 ;
        RECT  0.100 1.860 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.260 -0.140 2.540 0.320 ;
        RECT  1.220 -0.140 1.420 0.640 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END NR3M4HM

MACRO NR3M2HM
    CLASS CORE ;
    FOREIGN NR3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.580 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.140 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 1.080 0.700 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 1.840 1.900 2.060 ;
        RECT  1.740 0.440 1.900 2.060 ;
        RECT  0.620 0.620 1.900 0.820 ;
        RECT  1.640 0.440 1.900 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.220 1.800 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.140 -0.140 0.340 0.840 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END NR3M2HM

MACRO NR3M1HM
    CLASS CORE ;
    FOREIGN NR3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.580 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.140 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 1.080 0.700 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.370  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 1.840 1.900 2.060 ;
        RECT  1.740 0.440 1.900 2.060 ;
        RECT  0.620 0.620 1.900 0.820 ;
        RECT  1.640 0.440 1.900 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.220 1.800 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.140 -0.140 0.340 0.840 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END NR3M1HM

MACRO NR3M16HM
    CLASS CORE ;
    FOREIGN NR3M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.954  LAYER ME1  ;
        ANTENNAGATEAREA 0.954  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.897  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.060 5.900 1.260 ;
        LAYER ME2 ;
        RECT  5.700 0.840 5.900 1.560 ;
        LAYER ME1 ;
        RECT  4.320 1.000 7.480 1.160 ;
        RECT  5.600 1.000 6.000 1.320 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.954  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.700 0.980 11.120 1.150 ;
        RECT  7.700 0.980 7.900 1.560 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.954  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.990 3.840 1.190 ;
        RECT  0.100 0.840 0.300 1.190 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.735  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.220 1.580 11.500 2.060 ;
        RECT  11.300 0.340 11.500 2.060 ;
        RECT  0.820 0.660 11.500 0.820 ;
        RECT  11.220 0.340 11.500 0.820 ;
        RECT  8.060 1.580 11.500 1.740 ;
        RECT  10.180 0.340 10.460 0.820 ;
        RECT  9.140 0.340 9.420 0.820 ;
        RECT  8.100 0.340 8.380 0.820 ;
        RECT  7.060 0.340 7.340 0.820 ;
        RECT  6.020 0.340 6.300 0.820 ;
        RECT  4.980 0.340 5.260 0.820 ;
        RECT  3.940 0.340 4.220 0.820 ;
        RECT  2.900 0.340 3.180 0.820 ;
        RECT  1.860 0.340 2.140 0.820 ;
        RECT  0.820 0.340 1.100 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  3.420 1.900 3.700 2.540 ;
        RECT  2.380 1.900 2.660 2.540 ;
        RECT  1.340 1.900 1.620 2.540 ;
        RECT  0.300 1.900 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.700 -0.140 10.980 0.500 ;
        RECT  9.660 -0.140 9.940 0.500 ;
        RECT  8.620 -0.140 8.900 0.500 ;
        RECT  7.580 -0.140 7.860 0.500 ;
        RECT  6.540 -0.140 6.820 0.500 ;
        RECT  5.500 -0.140 5.780 0.500 ;
        RECT  4.460 -0.140 4.740 0.500 ;
        RECT  3.420 -0.140 3.700 0.500 ;
        RECT  2.380 -0.140 2.660 0.500 ;
        RECT  1.340 -0.140 1.620 0.500 ;
        RECT  0.300 -0.140 0.580 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.780 1.580 7.380 1.740 ;
        RECT  4.420 1.900 11.020 2.060 ;
        LAYER VTPH ;
        RECT  0.700 1.010 11.100 2.400 ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.010 ;
        RECT  0.000 0.000 0.700 1.140 ;
        RECT  11.100 0.000 11.600 1.140 ;
    END
END NR3M16HM

MACRO NR3M12HM
    CLASS CORE ;
    FOREIGN NR3M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.715  LAYER ME2  ;
        ANTENNAGATEAREA 0.715  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.352  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.040 4.700 1.240 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.360 ;
        LAYER ME1 ;
        RECT  3.480 0.980 4.960 1.360 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.715  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.700 0.980 7.900 1.560 ;
        RECT  7.220 0.980 7.900 1.260 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.715  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 1.300 1.260 ;
        RECT  0.100 0.840 0.300 1.260 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.092  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.020 1.740 8.300 2.060 ;
        RECT  8.100 0.340 8.300 2.060 ;
        RECT  0.740 0.660 8.300 0.820 ;
        RECT  8.020 0.340 8.300 0.820 ;
        RECT  5.940 1.580 7.300 1.740 ;
        RECT  6.980 0.340 7.260 0.820 ;
        RECT  5.940 0.340 6.220 1.740 ;
        RECT  4.900 0.340 5.180 0.820 ;
        RECT  3.860 0.340 4.140 0.820 ;
        RECT  2.820 0.340 3.100 0.820 ;
        RECT  1.780 0.340 2.060 0.820 ;
        RECT  0.740 0.340 1.020 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  2.300 1.900 2.580 2.540 ;
        RECT  1.260 1.900 1.540 2.540 ;
        RECT  0.220 1.900 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.500 -0.140 7.780 0.500 ;
        RECT  6.460 -0.140 6.740 0.500 ;
        RECT  5.420 -0.140 5.700 0.500 ;
        RECT  4.380 -0.140 4.660 0.500 ;
        RECT  3.340 -0.140 3.620 0.500 ;
        RECT  2.300 -0.140 2.580 0.500 ;
        RECT  1.260 -0.140 1.540 0.500 ;
        RECT  0.220 -0.140 0.500 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.700 1.580 5.220 1.740 ;
        RECT  3.300 1.900 7.820 2.060 ;
        LAYER VTPH ;
        RECT  0.580 0.960 7.940 2.400 ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 0.960 ;
        RECT  0.000 0.000 0.580 1.140 ;
        RECT  7.940 0.000 8.400 1.140 ;
    END
END NR3M12HM

MACRO NR3M0HM
    CLASS CORE ;
    FOREIGN NR3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.580 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.140 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 1.080 0.700 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.336  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 1.840 1.900 2.060 ;
        RECT  1.740 0.440 1.900 2.060 ;
        RECT  0.620 0.620 1.900 0.820 ;
        RECT  1.640 0.440 1.900 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.220 1.800 0.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.140 -0.140 0.340 0.840 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END NR3M0HM

MACRO NR3B1M8HM
    CLASS CORE ;
    FOREIGN NR3B1M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.476  LAYER ME2  ;
        ANTENNAGATEAREA 0.476  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.965  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.100 5.900 1.300 ;
        LAYER ME2 ;
        RECT  5.700 1.040 5.900 1.560 ;
        LAYER ME1 ;
        RECT  5.140 1.040 6.620 1.360 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.476  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.260 4.840 1.420 ;
        RECT  4.520 1.080 4.840 1.420 ;
        RECT  2.600 1.120 3.240 1.420 ;
        RECT  2.840 1.120 3.100 1.560 ;
        RECT  1.140 1.020 1.380 1.420 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.220 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.294  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.180 1.580 7.100 1.740 ;
        RECT  6.900 0.660 7.100 1.740 ;
        RECT  5.220 0.660 7.100 0.820 ;
        RECT  6.260 0.300 6.540 0.820 ;
        RECT  5.220 0.300 5.500 0.820 ;
        RECT  1.860 0.480 5.500 0.640 ;
        RECT  3.860 0.300 4.140 0.640 ;
        RECT  2.740 0.310 3.020 0.640 ;
        RECT  1.620 0.300 2.020 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  3.620 1.900 3.900 2.540 ;
        RECT  1.940 1.900 2.220 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.780 -0.140 7.060 0.500 ;
        RECT  5.740 -0.140 6.020 0.500 ;
        RECT  4.420 -0.140 4.700 0.320 ;
        RECT  3.300 -0.140 3.580 0.320 ;
        RECT  2.180 -0.140 2.460 0.320 ;
        RECT  1.100 -0.140 1.380 0.500 ;
        RECT  0.140 -0.140 0.340 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.380 0.900 0.660 ;
        RECT  0.740 0.700 1.700 0.860 ;
        RECT  1.540 0.800 4.080 0.960 ;
        RECT  3.440 0.800 4.080 1.080 ;
        RECT  0.740 0.380 0.900 2.060 ;
        RECT  0.620 1.540 0.900 2.060 ;
        RECT  1.100 1.580 2.580 1.740 ;
        RECT  3.260 1.580 4.980 1.740 ;
        RECT  1.100 1.580 1.380 1.800 ;
        RECT  2.420 1.720 3.420 1.880 ;
        RECT  4.700 1.580 4.980 2.060 ;
        RECT  4.700 1.900 7.100 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END NR3B1M8HM

MACRO NR3B1M4HM
    CLASS CORE ;
    FOREIGN NR3B1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.009  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.140 2.300 1.340 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.000 1.120 2.640 1.370 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.800 1.120 3.120 1.320 ;
        RECT  1.640 1.580 3.000 1.740 ;
        RECT  2.800 1.120 3.000 1.740 ;
        RECT  1.640 1.580 1.960 1.900 ;
        RECT  1.640 1.120 1.840 1.900 ;
        RECT  1.520 1.120 1.840 1.320 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.900 0.800 1.400 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.686  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.160 1.580 3.900 1.740 ;
        RECT  3.700 0.420 3.900 1.740 ;
        RECT  2.460 0.480 3.900 0.640 ;
        RECT  3.620 0.420 3.900 0.640 ;
        RECT  2.140 1.900 3.320 2.060 ;
        RECT  3.160 1.580 3.320 2.060 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  2.020 -0.140 2.220 0.640 ;
        RECT  0.380 -0.140 0.580 0.730 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.540 1.900 3.820 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.860 0.490 1.280 0.690 ;
        RECT  1.080 0.800 3.540 0.960 ;
        RECT  3.380 0.800 3.540 1.360 ;
        RECT  1.080 0.490 1.280 1.740 ;
        RECT  0.340 1.580 1.280 1.740 ;
        RECT  0.340 1.580 0.620 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END NR3B1M4HM

MACRO NR3B1M2HM
    CLASS CORE ;
    FOREIGN NR3B1M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.040 1.900 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.040 2.300 1.560 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 0.840 1.400 ;
        RECT  0.100 1.080 0.300 1.560 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.900 2.700 2.060 ;
        RECT  2.500 0.300 2.700 2.060 ;
        RECT  1.540 0.680 2.700 0.880 ;
        RECT  2.480 0.300 2.700 0.880 ;
        RECT  1.540 0.320 1.740 0.880 ;
        RECT  1.380 0.320 1.740 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.520 ;
        RECT  0.860 -0.140 1.140 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.300 0.300 0.500 0.880 ;
        RECT  0.300 0.680 1.360 0.880 ;
        RECT  0.620 1.580 1.360 1.740 ;
        RECT  1.160 0.680 1.360 1.740 ;
        RECT  0.340 1.720 0.780 1.940 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END NR3B1M2HM

MACRO NR3B1M1HM
    CLASS CORE ;
    FOREIGN NR3B1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.000 1.900 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.000 2.300 1.560 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.780 1.320 ;
        RECT  0.100 1.040 0.300 1.560 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.412  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.900 2.700 2.060 ;
        RECT  2.500 0.530 2.700 2.060 ;
        RECT  1.340 0.680 2.700 0.840 ;
        RECT  2.480 0.530 2.700 0.840 ;
        RECT  1.340 0.540 1.540 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.820 -0.140 2.100 0.320 ;
        RECT  0.700 -0.140 0.980 0.340 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 0.540 0.420 0.880 ;
        RECT  0.220 0.680 1.160 0.880 ;
        RECT  0.960 1.220 1.380 1.420 ;
        RECT  0.560 1.580 1.160 1.740 ;
        RECT  0.960 0.680 1.160 1.740 ;
        RECT  0.300 1.720 0.720 1.880 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.180 2.400 ;
        RECT  2.300 1.140 2.800 2.400 ;
        RECT  0.000 1.180 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
        RECT  1.180 0.000 2.300 1.180 ;
    END
END NR3B1M1HM

MACRO NR3B1M0HM
    CLASS CORE ;
    FOREIGN NR3B1M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.000 1.900 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.000 2.300 1.560 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.780 1.320 ;
        RECT  0.100 1.040 0.300 1.560 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.352  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.900 2.700 2.060 ;
        RECT  2.500 0.530 2.700 2.060 ;
        RECT  1.340 0.680 2.700 0.840 ;
        RECT  2.480 0.530 2.700 0.840 ;
        RECT  1.340 0.540 1.540 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.860 -0.140 2.060 0.380 ;
        RECT  0.820 -0.140 1.020 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 0.540 0.420 0.880 ;
        RECT  0.220 0.680 1.160 0.880 ;
        RECT  0.960 1.220 1.380 1.420 ;
        RECT  0.960 0.680 1.160 1.740 ;
        RECT  0.560 1.580 1.160 1.740 ;
        RECT  0.560 1.580 0.720 1.960 ;
        RECT  0.300 1.800 0.720 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END NR3B1M0HM

MACRO NR2M8HM
    CLASS CORE ;
    FOREIGN NR2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.080 2.800 1.280 ;
        RECT  2.100 0.800 2.300 1.280 ;
        RECT  0.800 0.800 2.300 0.960 ;
        RECT  0.800 0.800 1.000 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.960 1.260 3.900 1.420 ;
        RECT  3.620 0.840 3.900 1.420 ;
        RECT  0.320 1.440 3.120 1.600 ;
        RECT  2.960 1.260 3.120 1.600 ;
        RECT  1.600 1.120 1.880 1.600 ;
        RECT  0.320 1.060 0.520 1.600 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.273  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.580 4.300 1.740 ;
        RECT  4.100 0.480 4.300 1.740 ;
        RECT  3.140 0.480 4.300 0.640 ;
        RECT  0.900 1.760 3.440 1.920 ;
        RECT  3.280 1.580 3.440 1.920 ;
        RECT  2.460 0.720 3.300 0.880 ;
        RECT  3.140 0.480 3.300 0.880 ;
        RECT  2.460 0.480 2.620 0.880 ;
        RECT  0.940 0.480 2.620 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.620 1.900 3.900 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.960 -0.140 4.240 0.320 ;
        RECT  2.780 -0.140 2.980 0.560 ;
        RECT  1.540 -0.140 1.820 0.320 ;
        RECT  0.500 -0.140 0.700 0.660 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END NR2M8HM

MACRO NR2M6HM
    CLASS CORE ;
    FOREIGN NR2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.378  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.260 2.700 1.420 ;
        RECT  2.500 0.840 2.700 1.420 ;
        RECT  0.800 1.120 1.080 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.365  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.600 0.800 2.240 1.100 ;
        RECT  0.100 0.800 2.240 0.960 ;
        RECT  0.100 0.800 0.560 1.340 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.925  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.580 3.100 1.740 ;
        RECT  2.900 0.480 3.100 1.740 ;
        RECT  1.100 0.480 3.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        RECT  1.700 -0.140 1.980 0.320 ;
        RECT  0.660 -0.140 0.860 0.640 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END NR2M6HM

MACRO NR2M5HM
    CLASS CORE ;
    FOREIGN NR2M5HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.319  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 1.260 2.700 1.420 ;
        RECT  2.500 0.840 2.700 1.420 ;
        RECT  0.800 1.120 1.080 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.319  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.600 0.800 2.240 1.100 ;
        RECT  0.100 0.800 2.240 0.960 ;
        RECT  0.100 0.800 0.560 1.340 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.801  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.940 1.580 3.100 1.740 ;
        RECT  2.900 0.480 3.100 1.740 ;
        RECT  2.620 1.580 2.900 2.060 ;
        RECT  1.100 0.480 3.100 0.640 ;
        RECT  0.940 1.580 1.220 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        RECT  1.700 -0.140 1.980 0.320 ;
        RECT  0.660 -0.140 0.860 0.640 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END NR2M5HM

MACRO NR2M4HM
    CLASS CORE ;
    FOREIGN NR2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.031  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.180 1.070 1.380 1.270 ;
        LAYER ME2 ;
        RECT  1.180 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.760 1.060 1.440 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 1.440 1.900 1.600 ;
        RECT  1.660 1.060 1.900 1.600 ;
        RECT  0.300 1.060 0.500 1.600 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.760 2.300 1.920 ;
        RECT  2.100 0.500 2.300 1.920 ;
        RECT  0.620 0.500 2.300 0.800 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        RECT  0.160 -0.140 0.320 0.750 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END NR2M4HM

MACRO NR2M3HM
    CLASS CORE ;
    FOREIGN NR2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.400 1.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 1.320 1.900 1.480 ;
        RECT  1.680 1.040 1.900 1.480 ;
        RECT  0.500 1.320 0.700 1.960 ;
        RECT  0.300 1.050 0.500 1.480 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.438  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.660 2.300 1.800 ;
        RECT  1.340 1.640 2.300 1.800 ;
        RECT  1.640 0.660 2.300 0.820 ;
        RECT  1.640 0.370 1.800 0.820 ;
        RECT  1.420 0.370 1.800 0.530 ;
        RECT  0.900 1.730 1.500 1.890 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.820 1.960 2.100 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.980 -0.140 2.260 0.500 ;
        RECT  0.940 -0.140 1.220 0.500 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END NR2M3HM

MACRO NR2M2HM
    CLASS CORE ;
    FOREIGN NR2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.120 1.640 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 1.040 0.700 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.406  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.980 1.900 1.500 2.060 ;
        RECT  1.300 0.680 1.500 2.060 ;
        RECT  0.700 0.680 1.500 0.880 ;
        RECT  0.700 0.330 0.900 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  0.140 1.900 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  1.180 -0.140 1.460 0.500 ;
        RECT  0.180 -0.140 0.380 0.600 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END NR2M2HM

MACRO NR2M1HM
    CLASS CORE ;
    FOREIGN NR2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.030 1.140 1.570 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.220 0.600 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.321  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.020 1.840 1.500 2.100 ;
        RECT  1.300 0.610 1.500 2.100 ;
        RECT  0.700 0.610 1.500 0.770 ;
        RECT  0.700 0.490 0.980 0.770 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  0.140 1.840 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.100 -0.140 0.380 0.770 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END NR2M1HM

MACRO NR2M16HM
    CLASS CORE ;
    FOREIGN NR2M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.994  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.240 6.600 1.400 ;
        RECT  6.320 1.120 6.600 1.400 ;
        RECT  4.200 1.120 4.840 1.400 ;
        RECT  2.880 1.120 3.160 1.400 ;
        RECT  0.760 1.120 1.400 1.400 ;
        RECT  0.760 1.120 1.160 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.994  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.860 0.800 7.100 1.360 ;
        RECT  0.200 0.800 7.100 0.960 ;
        RECT  5.040 0.800 5.680 1.080 ;
        RECT  3.360 0.800 3.640 1.080 ;
        RECT  1.600 0.800 2.240 1.080 ;
        RECT  0.200 0.800 0.480 1.340 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.333  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.460 1.560 7.500 1.720 ;
        RECT  7.300 0.480 7.500 1.720 ;
        RECT  0.820 0.480 7.500 0.640 ;
        RECT  0.900 1.840 1.620 2.100 ;
        RECT  1.460 1.560 1.620 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.980 1.900 7.260 2.540 ;
        RECT  5.220 1.900 5.500 2.540 ;
        RECT  3.540 1.900 3.820 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.100 1.510 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.020 -0.140 7.300 0.320 ;
        RECT  5.900 -0.140 6.180 0.320 ;
        RECT  4.780 -0.140 5.060 0.320 ;
        RECT  3.660 -0.140 3.940 0.320 ;
        RECT  2.540 -0.140 2.820 0.320 ;
        RECT  1.420 -0.140 1.700 0.320 ;
        RECT  0.340 -0.140 0.620 0.640 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END NR2M16HM

MACRO NR2M12HM
    CLASS CORE ;
    FOREIGN NR2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.756  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.440 5.120 1.600 ;
        RECT  4.800 1.120 5.120 1.600 ;
        RECT  2.650 1.120 3.290 1.600 ;
        RECT  0.860 1.120 1.140 1.600 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.756  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.300 0.800 5.540 1.360 ;
        RECT  0.280 0.800 5.540 0.960 ;
        RECT  3.570 0.800 4.210 1.280 ;
        RECT  1.700 0.800 1.980 1.280 ;
        RECT  0.280 0.800 0.560 1.340 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.029  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.000 1.760 5.900 1.920 ;
        RECT  5.700 0.480 5.900 1.920 ;
        RECT  1.170 0.480 5.900 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.540 2.080 5.820 2.540 ;
        RECT  3.710 2.080 3.990 2.540 ;
        RECT  1.950 2.080 2.230 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.540 -0.140 5.820 0.320 ;
        RECT  4.420 -0.140 4.700 0.320 ;
        RECT  3.300 -0.140 3.580 0.320 ;
        RECT  2.180 -0.140 2.460 0.320 ;
        RECT  0.480 -0.140 0.760 0.320 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END NR2M12HM

MACRO NR2M0HM
    CLASS CORE ;
    FOREIGN NR2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.140 1.140 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.240 0.540 1.560 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.263  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.020 1.840 1.500 2.100 ;
        RECT  1.300 0.550 1.500 2.100 ;
        RECT  0.700 0.550 1.500 0.770 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  0.140 1.840 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.100 -0.140 0.380 0.770 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END NR2M0HM

MACRO NR2B1M8HM
    CLASS CORE ;
    FOREIGN NR2B1M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.080 0.800 3.800 1.100 ;
        RECT  1.400 0.800 3.800 0.960 ;
        RECT  1.400 0.800 1.620 1.280 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.900 0.760 1.280 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.580 4.700 1.740 ;
        RECT  4.500 0.480 4.700 1.740 ;
        RECT  1.580 0.480 4.700 0.640 ;
        RECT  1.580 1.900 2.260 2.100 ;
        RECT  2.100 1.580 2.260 2.100 ;
        RECT  1.580 0.300 1.860 0.640 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.420 -0.140 4.700 0.320 ;
        RECT  3.300 -0.140 3.580 0.320 ;
        RECT  2.180 -0.140 2.460 0.320 ;
        RECT  0.780 -0.140 1.060 0.320 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.360 1.900 4.640 2.540 ;
        RECT  2.420 1.900 2.700 2.540 ;
        RECT  0.740 1.900 1.020 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.220 0.530 1.140 0.740 ;
        RECT  1.780 1.120 2.880 1.420 ;
        RECT  4.020 1.060 4.300 1.420 ;
        RECT  1.780 1.260 4.300 1.420 ;
        RECT  0.980 0.530 1.140 1.740 ;
        RECT  0.220 1.540 1.140 1.740 ;
        RECT  1.780 1.120 1.940 1.740 ;
        RECT  0.220 1.550 1.940 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END NR2B1M8HM

MACRO NR2B1M4HM
    CLASS CORE ;
    FOREIGN NR2B1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.520 0.900 1.960 1.220 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.390 1.010 0.700 1.560 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.568  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.760 3.100 1.920 ;
        RECT  2.900 0.740 3.100 1.920 ;
        RECT  2.300 0.740 3.100 0.900 ;
        RECT  2.300 0.300 2.580 0.900 ;
        RECT  1.400 0.500 2.580 0.700 ;
        RECT  1.180 0.300 1.580 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.720 2.080 3.000 2.540 ;
        RECT  0.780 2.080 1.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.550 ;
        RECT  1.740 -0.140 2.020 0.320 ;
        RECT  0.660 -0.140 0.940 0.530 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.850 ;
        RECT  0.100 0.690 1.200 0.850 ;
        RECT  2.460 1.060 2.740 1.600 ;
        RECT  0.980 1.440 2.740 1.600 ;
        RECT  0.980 0.690 1.200 1.920 ;
        RECT  0.220 1.760 1.200 1.920 ;
        RECT  0.220 1.760 0.500 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END NR2B1M4HM

MACRO NR2B1M2HM
    CLASS CORE ;
    FOREIGN NR2B1M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.570 1.560 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.320 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.385  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.730 1.900 2.020 ;
        RECT  1.740 0.500 1.900 2.020 ;
        RECT  1.180 0.500 1.900 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.630 2.040 0.910 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.600 -0.140 0.890 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.020 0.680 ;
        RECT  0.820 0.480 1.020 1.720 ;
        RECT  0.100 1.520 1.020 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END NR2B1M2HM

MACRO NR2B1M1HM
    CLASS CORE ;
    FOREIGN NR2B1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.570 1.560 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.320 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.342  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.730 1.900 2.020 ;
        RECT  1.740 0.500 1.900 2.020 ;
        RECT  1.180 0.500 1.900 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.630 2.040 0.910 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.600 -0.140 0.890 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.020 0.680 ;
        RECT  0.820 0.480 1.020 1.720 ;
        RECT  0.100 1.520 1.020 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END NR2B1M1HM

MACRO NR2B1M12HM
    CLASS CORE ;
    FOREIGN NR2B1M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.744  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.800 1.260 5.760 1.420 ;
        RECT  5.480 1.120 5.760 1.420 ;
        RECT  3.580 1.120 3.860 1.420 ;
        RECT  1.800 1.260 2.360 1.560 ;
        RECT  1.800 0.980 2.080 1.560 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.256  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 1.080 1.360 ;
        RECT  0.100 1.040 0.400 1.560 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.664  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.520 1.580 6.700 1.740 ;
        RECT  6.500 0.480 6.700 1.740 ;
        RECT  2.650 0.480 6.700 0.640 ;
        RECT  2.410 0.300 2.810 0.500 ;
        RECT  1.980 1.820 2.680 2.100 ;
        RECT  2.520 1.580 2.680 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.300 1.900 6.580 2.540 ;
        RECT  4.520 1.900 4.800 2.540 ;
        RECT  2.840 1.900 3.120 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.840 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.340 -0.140 6.620 0.320 ;
        RECT  5.220 -0.140 5.500 0.320 ;
        RECT  4.100 -0.140 4.380 0.320 ;
        RECT  2.970 -0.140 3.250 0.320 ;
        RECT  1.890 -0.140 2.170 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.100 -0.140 0.380 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.360 0.900 0.820 ;
        RECT  0.620 0.660 2.480 0.820 ;
        RECT  2.310 0.800 6.340 0.960 ;
        RECT  2.310 0.800 3.060 1.100 ;
        RECT  4.340 0.800 4.620 1.100 ;
        RECT  6.120 0.800 6.340 1.300 ;
        RECT  1.360 0.660 1.560 1.740 ;
        RECT  0.620 1.580 1.560 1.740 ;
        RECT  0.620 1.580 0.900 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END NR2B1M12HM

MACRO NR2B1M0HM
    CLASS CORE ;
    FOREIGN NR2B1M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.040 1.570 1.560 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.320 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 1.730 1.900 2.020 ;
        RECT  1.740 0.500 1.900 2.020 ;
        RECT  1.180 0.500 1.900 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.630 2.040 0.910 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.600 -0.140 0.890 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.020 0.680 ;
        RECT  0.820 0.480 1.020 1.720 ;
        RECT  0.100 1.520 1.020 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END NR2B1M0HM

MACRO ND4M8HM
    CLASS CORE ;
    FOREIGN ND4M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.438  LAYER ME2  ;
        ANTENNAGATEAREA 0.438  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.508  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.150 3.100 1.350 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.480 1.150 3.480 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.438  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.680 1.120 7.160 1.560 ;
        RECT  6.040 1.120 7.160 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.438  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.640 1.150 5.040 1.350 ;
        RECT  3.640 0.840 3.960 1.350 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.438  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.150 1.960 1.420 ;
        RECT  0.440 1.150 0.760 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.764  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.660 0.790 7.020 0.950 ;
        RECT  6.740 0.540 7.020 0.950 ;
        RECT  6.260 1.580 6.460 1.990 ;
        RECT  1.060 1.580 6.460 1.740 ;
        RECT  5.660 0.620 5.980 0.950 ;
        RECT  5.660 0.620 5.880 1.740 ;
        RECT  5.220 1.580 5.420 1.990 ;
        RECT  4.180 1.580 4.380 1.990 ;
        RECT  3.140 1.580 3.340 1.990 ;
        RECT  2.100 1.580 2.300 1.990 ;
        RECT  1.060 1.580 1.260 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.740 1.900 7.020 2.540 ;
        RECT  5.700 1.900 5.980 2.540 ;
        RECT  4.660 1.900 4.940 2.540 ;
        RECT  3.620 1.900 3.900 2.540 ;
        RECT  2.580 1.900 2.860 2.540 ;
        RECT  1.540 1.900 1.820 2.540 ;
        RECT  0.540 1.730 0.740 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  1.540 -0.140 1.820 0.500 ;
        RECT  0.500 -0.140 0.780 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.060 0.300 1.260 0.990 ;
        RECT  2.100 0.300 2.300 0.990 ;
        RECT  3.100 0.620 3.380 0.990 ;
        RECT  1.060 0.830 3.380 0.990 ;
        RECT  2.580 0.300 4.940 0.460 ;
        RECT  2.580 0.300 2.860 0.500 ;
        RECT  3.620 0.300 3.900 0.500 ;
        RECT  4.660 0.300 4.940 0.500 ;
        RECT  5.180 0.300 6.500 0.460 ;
        RECT  6.220 0.300 6.500 0.630 ;
        RECT  4.140 0.620 4.420 0.940 ;
        RECT  5.180 0.300 5.420 0.940 ;
        RECT  4.140 0.780 5.420 0.940 ;
        LAYER VTPH ;
        RECT  0.000 1.280 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.280 ;
    END
END ND4M8HM

MACRO ND4M6HM
    CLASS CORE ;
    FOREIGN ND4M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        ANTENNAGATEAREA 0.071  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.508  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.820 1.080 2.020 1.280 ;
        LAYER ME2 ;
        RECT  1.700 0.980 2.020 1.560 ;
        LAYER ME1 ;
        RECT  1.820 0.980 2.090 1.460 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        ANTENNAGATEAREA 0.071  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.582  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.800 0.940 1.000 1.140 ;
        LAYER ME2 ;
        RECT  0.800 0.800 1.100 1.390 ;
        LAYER ME1 ;
        RECT  0.780 0.830 1.020 1.350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.600 1.160 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.660 0.460 5.900 2.100 ;
        RECT  4.620 1.460 5.900 1.660 ;
        RECT  4.580 0.660 5.900 0.860 ;
        RECT  5.620 0.460 5.900 0.860 ;
        RECT  4.580 0.470 4.860 0.860 ;
        RECT  4.620 1.460 4.820 2.100 ;
        END
    END Z
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        ANTENNAGATEAREA 0.071  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.362  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.080 2.570 1.280 ;
        LAYER ME2 ;
        RECT  2.370 0.800 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.250 0.980 2.570 1.390 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.100 1.880 5.380 2.540 ;
        RECT  4.100 1.460 4.300 2.540 ;
        RECT  0.100 1.630 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.380 0.500 ;
        RECT  4.060 -0.140 4.340 0.690 ;
        RECT  3.590 -0.140 3.870 0.500 ;
        RECT  2.470 -0.140 2.750 0.500 ;
        RECT  0.140 -0.140 0.420 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.500 0.300 1.760 0.820 ;
        RECT  1.500 0.660 2.950 0.820 ;
        RECT  2.730 0.660 2.950 1.260 ;
        RECT  1.500 0.300 1.660 1.780 ;
        RECT  1.500 1.620 2.220 1.780 ;
        RECT  1.020 0.300 1.340 0.560 ;
        RECT  3.170 1.040 3.490 1.240 ;
        RECT  0.660 1.640 1.340 1.800 ;
        RECT  1.180 0.300 1.340 2.100 ;
        RECT  3.170 1.040 3.330 2.100 ;
        RECT  1.180 1.940 3.330 2.100 ;
        RECT  3.110 0.350 3.310 0.820 ;
        RECT  3.110 0.660 3.870 0.820 ;
        RECT  3.710 1.050 5.460 1.210 ;
        RECT  3.710 0.660 3.870 2.100 ;
        RECT  3.490 1.460 3.870 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END ND4M6HM

MACRO ND4M4HM
    CLASS CORE ;
    FOREIGN ND4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        ANTENNAGATEAREA 0.228  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.075  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.150 1.900 1.350 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.480 1.150 2.120 1.420 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        ANTENNAGATEAREA 0.228  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.144  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.150 3.100 1.350 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.800 1.150 3.540 1.350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.860 1.120 5.100 1.560 ;
        RECT  4.480 1.120 5.100 1.420 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.150 1.080 1.420 ;
        RECT  0.100 1.150 0.360 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.220 1.580 4.500 2.100 ;
        RECT  4.160 0.620 4.500 0.840 ;
        RECT  4.160 0.620 4.320 1.740 ;
        RECT  0.620 1.580 4.500 1.740 ;
        RECT  3.180 1.580 3.460 2.100 ;
        RECT  1.660 1.580 1.940 2.100 ;
        RECT  0.620 1.580 0.900 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.740 1.900 5.020 2.540 ;
        RECT  3.700 1.900 3.980 2.540 ;
        RECT  2.650 1.900 2.930 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.820 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.620 0.380 0.840 ;
        RECT  1.140 0.620 1.420 0.840 ;
        RECT  0.100 0.660 1.420 0.840 ;
        RECT  2.180 0.620 2.460 0.840 ;
        RECT  0.100 0.680 2.460 0.840 ;
        RECT  1.660 0.300 3.460 0.460 ;
        RECT  1.660 0.300 1.940 0.520 ;
        RECT  3.180 0.300 3.460 0.520 ;
        RECT  3.700 0.300 5.100 0.460 ;
        RECT  4.820 0.300 5.100 0.520 ;
        RECT  2.660 0.620 2.940 0.840 ;
        RECT  3.700 0.300 3.980 0.840 ;
        RECT  2.660 0.680 3.980 0.840 ;
        LAYER VTPH ;
        RECT  0.000 1.280 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.280 ;
    END
END ND4M4HM

MACRO ND4M2HM
    CLASS CORE ;
    FOREIGN ND4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 1.130 2.300 1.350 ;
        RECT  2.080 0.840 2.300 1.350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.600 1.350 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.350 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.130 0.560 1.410 ;
        RECT  0.100 1.130 0.360 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.502  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.620 1.580 2.700 1.740 ;
        RECT  2.500 0.300 2.700 1.740 ;
        RECT  2.180 0.300 2.700 0.660 ;
        RECT  1.660 1.580 1.940 2.100 ;
        RECT  0.620 1.580 0.900 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.730 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.100 -0.140 0.380 0.670 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND4M2HM

MACRO ND4M1HM
    CLASS CORE ;
    FOREIGN ND4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.810 2.320 1.270 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.810 1.720 1.270 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.810 1.100 1.270 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.810 0.560 1.270 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.397  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.490 2.700 1.740 ;
        RECT  2.500 0.300 2.700 1.740 ;
        RECT  2.180 0.300 2.700 0.550 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.380 2.020 2.660 2.540 ;
        RECT  1.220 2.020 1.500 2.540 ;
        RECT  0.100 2.020 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.100 -0.140 0.380 0.500 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND4M1HM

MACRO ND4M16HM
    CLASS CORE ;
    FOREIGN ND4M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.887  LAYER ME1  ;
        ANTENNAGATEAREA 0.887  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.589  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.160 4.700 1.360 ;
        LAYER ME2 ;
        RECT  4.500 1.040 4.700 1.560 ;
        LAYER ME1 ;
        RECT  3.700 1.150 6.140 1.420 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.887  LAYER ME1  ;
        ANTENNAGATEAREA 0.887  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.589  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.160 8.300 1.360 ;
        LAYER ME2 ;
        RECT  8.100 1.040 8.300 1.560 ;
        LAYER ME1 ;
        RECT  7.300 1.150 9.740 1.420 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.865  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.200 1.120 13.500 1.560 ;
        RECT  11.130 1.120 13.500 1.420 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.865  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.150 3.020 1.420 ;
        RECT  0.100 1.150 0.360 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.356  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.420 0.690 12.820 0.910 ;
        RECT  12.580 1.580 12.780 1.990 ;
        RECT  0.660 1.580 12.780 1.740 ;
        RECT  11.540 1.580 11.740 1.990 ;
        RECT  10.500 0.690 10.700 1.990 ;
        RECT  10.420 0.690 10.700 1.740 ;
        RECT  9.460 1.580 9.660 1.990 ;
        RECT  8.420 1.580 8.620 1.990 ;
        RECT  7.380 1.580 7.580 1.990 ;
        RECT  5.860 1.580 6.060 1.990 ;
        RECT  4.820 1.580 5.020 1.990 ;
        RECT  3.780 1.580 3.980 1.990 ;
        RECT  2.740 1.580 2.940 1.990 ;
        RECT  1.700 1.580 1.900 1.990 ;
        RECT  0.660 1.580 0.860 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  13.060 1.900 13.340 2.540 ;
        RECT  12.020 1.900 12.300 2.540 ;
        RECT  10.980 1.900 11.260 2.540 ;
        RECT  9.940 1.900 10.220 2.540 ;
        RECT  8.900 1.900 9.180 2.540 ;
        RECT  7.860 1.900 8.140 2.540 ;
        RECT  6.340 1.900 6.980 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.730 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.410 0.340 0.920 ;
        RECT  1.180 0.340 1.380 0.920 ;
        RECT  2.220 0.320 2.420 0.920 ;
        RECT  3.260 0.320 3.460 0.920 ;
        RECT  0.140 0.710 6.620 0.920 ;
        RECT  3.700 0.320 9.740 0.500 ;
        RECT  9.940 0.320 13.380 0.530 ;
        RECT  9.940 0.320 10.220 0.990 ;
        RECT  6.820 0.760 10.220 0.990 ;
        LAYER VTPH ;
        RECT  1.660 1.280 5.080 2.400 ;
        RECT  8.370 1.280 11.780 2.400 ;
        RECT  0.000 1.320 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.280 ;
        RECT  0.000 0.000 1.660 1.320 ;
        RECT  5.080 0.000 8.370 1.320 ;
        RECT  11.780 0.000 13.600 1.320 ;
    END
END ND4M16HM

MACRO ND4M12HM
    CLASS CORE ;
    FOREIGN ND4M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.683  LAYER ME1  ;
        ANTENNAGATEAREA 0.683  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.523  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.150 4.300 1.350 ;
        LAYER ME2 ;
        RECT  4.100 1.040 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.160 1.150 4.890 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.683  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.440 1.120 10.760 1.560 ;
        RECT  9.070 1.120 10.760 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.683  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.240 1.150 7.860 1.420 ;
        RECT  5.240 0.840 5.560 1.420 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.683  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.150 2.660 1.420 ;
        RECT  0.100 1.150 0.360 1.560 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.609  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.420 0.660 10.780 0.820 ;
        RECT  10.500 0.520 10.780 0.820 ;
        RECT  10.020 1.580 10.220 1.990 ;
        RECT  0.660 1.580 10.220 1.740 ;
        RECT  8.980 1.580 9.180 1.990 ;
        RECT  8.420 0.660 8.760 1.740 ;
        RECT  7.940 1.580 8.140 1.990 ;
        RECT  6.900 1.580 7.100 1.990 ;
        RECT  5.860 1.580 6.060 1.990 ;
        RECT  4.820 1.580 5.020 1.990 ;
        RECT  3.780 1.580 3.980 1.990 ;
        RECT  2.740 1.580 2.940 1.990 ;
        RECT  1.700 1.580 1.900 1.990 ;
        RECT  0.660 1.580 0.860 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.500 1.900 10.780 2.540 ;
        RECT  9.460 1.900 9.740 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.730 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.100 -0.140 0.380 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.470 0.860 0.920 ;
        RECT  0.660 0.700 5.060 0.920 ;
        RECT  3.180 0.320 7.700 0.500 ;
        RECT  7.900 0.320 10.300 0.500 ;
        RECT  7.900 0.320 8.180 0.960 ;
        RECT  5.820 0.740 8.180 0.960 ;
        LAYER VTPH ;
        RECT  0.000 1.290 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.290 ;
    END
END ND4M12HM

MACRO ND4M0HM
    CLASS CORE ;
    FOREIGN ND4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.840 2.320 1.270 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.660 1.330 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.100 1.330 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.330 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.346  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.490 2.700 1.740 ;
        RECT  2.500 0.300 2.700 1.740 ;
        RECT  2.180 0.300 2.700 0.550 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.380 2.020 2.660 2.540 ;
        RECT  1.220 2.020 1.500 2.540 ;
        RECT  0.100 2.020 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.100 -0.140 0.380 0.500 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND4M0HM

MACRO ND4B2M8HM
    CLASS CORE ;
    FOREIGN ND4B2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER ME1  ;
        ANTENNAGATEAREA 0.445  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.495  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.180 5.100 1.380 ;
        LAYER ME2 ;
        RECT  4.900 1.040 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.660 1.140 5.660 1.420 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER ME1  ;
        ANTENNAGATEAREA 0.445  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.495  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.180 3.900 1.380 ;
        LAYER ME2 ;
        RECT  3.700 1.040 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.100 1.140 4.100 1.420 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 0.500 1.560 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.120 1.040 8.700 1.560 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.736  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 0.660 7.630 0.860 ;
        RECT  7.360 0.470 7.630 0.860 ;
        RECT  6.880 1.580 7.080 1.990 ;
        RECT  1.680 1.580 7.080 1.740 ;
        RECT  6.100 0.660 6.300 1.740 ;
        RECT  5.840 1.580 6.040 1.990 ;
        RECT  4.800 1.580 5.000 1.990 ;
        RECT  3.760 1.580 3.960 1.990 ;
        RECT  2.720 1.580 2.920 1.990 ;
        RECT  1.680 1.580 1.880 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.360 1.900 7.640 2.540 ;
        RECT  6.320 1.900 6.600 2.540 ;
        RECT  5.280 1.900 5.560 2.540 ;
        RECT  4.240 1.900 4.520 2.540 ;
        RECT  3.200 1.900 3.480 2.540 ;
        RECT  2.160 1.900 2.440 2.540 ;
        RECT  1.120 1.900 1.400 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.380 -0.140 8.620 0.680 ;
        RECT  2.160 -0.140 2.440 0.500 ;
        RECT  1.120 -0.140 1.400 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.410 0.380 0.820 ;
        RECT  0.100 0.660 0.920 0.820 ;
        RECT  0.720 1.140 2.540 1.420 ;
        RECT  0.720 0.660 0.920 2.100 ;
        RECT  0.100 1.820 0.920 2.100 ;
        RECT  1.640 0.720 4.000 0.940 ;
        RECT  3.200 0.300 5.560 0.500 ;
        RECT  4.240 0.300 4.520 0.860 ;
        RECT  5.740 0.300 7.120 0.500 ;
        RECT  5.740 0.300 5.940 0.940 ;
        RECT  4.760 0.740 5.940 0.940 ;
        RECT  7.800 0.410 8.140 0.690 ;
        RECT  6.620 1.140 7.960 1.420 ;
        RECT  7.800 0.410 7.960 2.060 ;
        RECT  7.800 1.860 8.660 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.030 2.400 ;
        RECT  7.730 1.140 8.800 2.400 ;
        RECT  0.000 1.300 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
        RECT  1.030 0.000 7.730 1.300 ;
    END
END ND4B2M8HM

MACRO ND4B2M4HM
    CLASS CORE ;
    FOREIGN ND4B2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.440 5.100 1.600 ;
        RECT  4.760 1.020 5.100 1.600 ;
        RECT  3.260 1.120 3.540 1.600 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.480 0.840 2.200 1.280 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.760 1.260 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.580 0.980 6.300 1.300 ;
        RECT  6.080 0.840 6.300 1.300 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.100 1.760 4.860 1.920 ;
        RECT  2.900 0.800 4.260 0.960 ;
        RECT  3.980 0.620 4.260 0.960 ;
        RECT  2.900 0.800 3.100 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.060 1.860 5.340 2.540 ;
        RECT  3.980 2.080 4.260 2.540 ;
        RECT  2.840 2.080 3.120 2.540 ;
        RECT  1.700 2.080 1.980 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.860 -0.140 6.140 0.560 ;
        RECT  2.620 -0.140 2.900 0.320 ;
        RECT  0.720 -0.140 1.000 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.640 ;
        RECT  0.100 0.480 1.220 0.640 ;
        RECT  1.020 0.480 1.220 1.600 ;
        RECT  2.420 1.100 2.700 1.600 ;
        RECT  0.140 1.440 2.700 1.600 ;
        RECT  0.140 1.440 0.340 2.060 ;
        RECT  3.100 0.300 5.140 0.460 ;
        RECT  1.700 0.300 1.980 0.640 ;
        RECT  4.860 0.300 5.140 0.500 ;
        RECT  3.100 0.300 3.380 0.640 ;
        RECT  1.700 0.480 3.380 0.640 ;
        RECT  5.340 0.300 5.620 0.820 ;
        RECT  4.440 0.660 5.620 0.820 ;
        RECT  4.440 0.660 4.600 1.280 ;
        RECT  3.720 1.120 4.600 1.280 ;
        RECT  5.260 0.660 5.420 1.620 ;
        RECT  5.260 1.460 5.860 1.620 ;
        RECT  5.580 1.460 5.860 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.370 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.370 ;
    END
END ND4B2M4HM

MACRO ND4B2M2HM
    CLASS CORE ;
    FOREIGN ND4B2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 0.820 2.300 1.220 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.820 1.720 1.220 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.300 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.400 1.080 3.900 1.560 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.502  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.340 2.900 0.500 ;
        RECT  2.260 1.580 2.700 2.060 ;
        RECT  2.500 0.340 2.700 2.060 ;
        RECT  1.420 1.580 2.700 1.740 ;
        RECT  1.180 1.900 1.580 2.060 ;
        RECT  1.420 1.580 1.580 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  1.740 1.900 2.020 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.340 0.380 ;
        RECT  0.720 -0.140 1.000 0.340 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.430 0.380 0.660 ;
        RECT  0.100 0.500 1.140 0.660 ;
        RECT  0.920 0.500 1.140 1.740 ;
        RECT  0.140 1.580 1.140 1.740 ;
        RECT  0.140 1.580 0.340 2.000 ;
        RECT  3.620 0.520 3.900 0.820 ;
        RECT  2.860 0.660 3.900 0.820 ;
        RECT  2.860 0.660 3.060 1.880 ;
        RECT  2.860 1.720 3.900 1.880 ;
        RECT  3.620 1.720 3.900 2.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END ND4B2M2HM

MACRO ND4B2M1HM
    CLASS CORE ;
    FOREIGN ND4B2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 0.790 2.300 1.350 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.790 1.720 1.220 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.300 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.620 0.840 3.900 1.370 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.431  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.340 2.900 0.560 ;
        RECT  2.480 1.660 2.740 2.100 ;
        RECT  2.500 0.340 2.740 2.100 ;
        RECT  1.300 1.660 2.740 1.920 ;
        RECT  1.300 1.660 1.560 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.260 2.080 3.900 2.540 ;
        RECT  1.880 2.080 2.160 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  0.720 -0.140 1.000 0.340 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.430 0.380 0.660 ;
        RECT  0.100 0.500 1.140 0.660 ;
        RECT  0.920 0.500 1.140 1.740 ;
        RECT  0.100 1.580 1.140 1.740 ;
        RECT  0.100 1.580 0.380 2.000 ;
        RECT  3.620 0.300 3.900 0.660 ;
        RECT  3.240 0.500 3.900 0.660 ;
        RECT  2.900 0.910 3.400 1.190 ;
        RECT  3.240 0.500 3.400 1.750 ;
        RECT  3.240 1.530 3.900 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END ND4B2M1HM

MACRO ND4B2M0HM
    CLASS CORE ;
    FOREIGN ND4B2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 0.800 2.300 1.320 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.810 1.720 1.220 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.300 ;
        END
    END NA
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.620 0.840 3.900 1.300 ;
        END
    END NB
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.380  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.340 2.900 0.560 ;
        RECT  2.500 0.340 2.740 2.100 ;
        RECT  1.320 1.660 2.740 1.830 ;
        RECT  1.320 1.660 1.580 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.260 2.080 3.900 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  0.720 -0.140 1.000 0.340 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.420 0.380 0.680 ;
        RECT  0.100 0.500 1.140 0.680 ;
        RECT  0.920 0.500 1.140 1.740 ;
        RECT  0.100 1.580 1.140 1.740 ;
        RECT  0.100 1.580 0.380 2.000 ;
        RECT  3.620 0.300 3.900 0.660 ;
        RECT  3.240 0.500 3.900 0.660 ;
        RECT  2.900 0.910 3.400 1.190 ;
        RECT  3.240 0.500 3.400 1.750 ;
        RECT  3.240 1.530 3.900 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END ND4B2M0HM

MACRO ND4B1M8HM
    CLASS CORE ;
    FOREIGN ND4B1M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER ME1  ;
        ANTENNAGATEAREA 0.445  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.495  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.150 3.900 1.350 ;
        LAYER ME2 ;
        RECT  3.700 1.040 3.900 1.560 ;
        LAYER ME1 ;
        RECT  3.100 1.110 4.100 1.390 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER ME1  ;
        ANTENNAGATEAREA 0.445  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.495  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 1.150 5.100 1.350 ;
        LAYER ME2 ;
        RECT  4.900 1.040 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.660 1.110 5.660 1.390 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 1.110 7.600 1.560 ;
        RECT  6.700 1.110 7.600 1.390 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.760 1.270 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.776  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.280 0.670 7.680 0.950 ;
        RECT  6.840 1.580 7.120 2.100 ;
        RECT  1.640 1.580 7.120 1.740 ;
        RECT  6.280 0.670 6.540 1.740 ;
        RECT  5.800 1.580 6.080 2.100 ;
        RECT  4.760 1.580 5.040 2.100 ;
        RECT  3.720 1.580 4.000 2.100 ;
        RECT  2.680 1.580 2.960 2.100 ;
        RECT  1.640 1.580 1.920 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.360 1.900 7.640 2.540 ;
        RECT  6.320 1.900 6.600 2.540 ;
        RECT  5.280 1.900 5.560 2.540 ;
        RECT  4.240 1.900 4.520 2.540 ;
        RECT  3.200 1.900 3.480 2.540 ;
        RECT  2.160 1.900 2.440 2.540 ;
        RECT  1.120 1.900 1.400 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  2.200 -0.140 2.480 0.500 ;
        RECT  0.620 -0.140 1.400 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.410 0.380 0.680 ;
        RECT  0.100 0.520 1.470 0.680 ;
        RECT  1.260 0.520 1.470 1.390 ;
        RECT  1.260 1.110 2.540 1.390 ;
        RECT  1.260 0.520 1.460 1.740 ;
        RECT  0.100 1.580 1.460 1.740 ;
        RECT  0.100 1.580 0.380 2.100 ;
        RECT  1.680 0.300 1.960 0.820 ;
        RECT  2.720 0.300 3.000 0.820 ;
        RECT  1.680 0.660 4.080 0.820 ;
        RECT  3.240 0.300 5.600 0.500 ;
        RECT  4.280 0.300 4.560 0.860 ;
        RECT  5.840 0.300 7.160 0.500 ;
        RECT  5.840 0.300 6.120 0.820 ;
        RECT  4.760 0.660 6.120 0.820 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.030 2.400 ;
        RECT  0.000 1.300 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
        RECT  1.030 0.000 8.400 1.300 ;
    END
END ND4B1M8HM

MACRO ND4B1M4HM
    CLASS CORE ;
    FOREIGN ND4B1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.480 1.000 2.200 1.280 ;
        RECT  1.480 0.840 1.960 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.050 4.040 1.330 ;
        RECT  3.300 1.050 3.500 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.160 1.050 5.500 1.560 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.800 0.760 1.280 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.848  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.620 0.620 4.900 1.920 ;
        RECT  3.720 1.550 4.900 1.710 ;
        RECT  4.500 0.620 4.900 1.710 ;
        RECT  1.100 1.760 3.900 1.920 ;
        RECT  3.720 1.550 3.900 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.140 1.870 5.420 2.540 ;
        RECT  4.100 1.870 4.380 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  1.700 2.080 1.980 2.540 ;
        RECT  0.620 1.870 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  2.580 -0.140 2.860 0.500 ;
        RECT  0.720 -0.140 1.000 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.640 ;
        RECT  0.100 0.480 1.220 0.640 ;
        RECT  1.020 0.480 1.220 1.600 ;
        RECT  2.420 1.050 2.700 1.600 ;
        RECT  0.140 1.440 2.700 1.600 ;
        RECT  0.140 1.440 0.340 2.060 ;
        RECT  1.700 0.340 2.420 0.620 ;
        RECT  2.260 0.340 2.420 0.820 ;
        RECT  3.580 0.620 3.860 0.820 ;
        RECT  2.260 0.660 3.860 0.820 ;
        RECT  3.060 0.300 5.420 0.460 ;
        RECT  3.060 0.300 3.340 0.500 ;
        RECT  4.100 0.300 4.380 0.500 ;
        RECT  5.140 0.300 5.420 0.500 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END ND4B1M4HM

MACRO ND4B1M2HM
    CLASS CORE ;
    FOREIGN ND4B1M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 0.810 1.900 1.270 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.080 0.810 2.340 1.260 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.750 2.720 1.260 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.410 0.830 0.760 1.290 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.525  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.580 3.100 1.740 ;
        RECT  2.900 0.300 3.100 1.740 ;
        RECT  2.680 0.300 3.100 0.520 ;
        RECT  2.300 1.580 2.570 2.060 ;
        RECT  1.260 1.580 1.530 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 1.900 3.100 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.740 1.900 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  0.840 -0.140 1.120 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 0.300 0.520 0.660 ;
        RECT  0.240 0.480 1.100 0.660 ;
        RECT  0.920 0.940 1.340 1.220 ;
        RECT  0.920 0.480 1.100 1.740 ;
        RECT  0.100 1.580 1.100 1.740 ;
        RECT  0.100 1.580 0.380 2.010 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END ND4B1M2HM

MACRO ND4B1M1HM
    CLASS CORE ;
    FOREIGN ND4B1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 0.770 1.900 1.270 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.080 0.770 2.300 1.260 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.770 2.720 1.260 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.370 0.830 0.760 1.160 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.497  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.680 3.100 1.840 ;
        RECT  2.900 0.300 3.100 1.840 ;
        RECT  2.680 0.300 3.100 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 2.080 3.100 2.540 ;
        RECT  1.710 2.080 1.990 2.540 ;
        RECT  0.580 2.080 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  0.840 -0.140 1.120 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 0.300 0.520 0.660 ;
        RECT  0.240 0.480 1.100 0.660 ;
        RECT  0.920 0.940 1.340 1.220 ;
        RECT  0.920 0.480 1.100 1.480 ;
        RECT  0.100 1.320 1.100 1.480 ;
        RECT  0.100 1.320 0.380 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END ND4B1M1HM

MACRO ND4B1M0HM
    CLASS CORE ;
    FOREIGN ND4B1M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 0.790 1.900 1.270 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.080 0.790 2.300 1.260 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.062  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.790 2.720 1.260 ;
        END
    END D
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.830 0.760 1.160 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 1.620 3.100 1.780 ;
        RECT  2.900 0.300 3.100 1.780 ;
        RECT  2.680 0.300 3.100 0.520 ;
        RECT  2.260 1.620 2.540 1.940 ;
        RECT  1.180 1.620 1.460 1.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 2.020 3.100 2.540 ;
        RECT  1.710 2.020 1.990 2.540 ;
        RECT  0.580 2.020 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  0.840 -0.140 1.120 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 0.300 0.520 0.660 ;
        RECT  0.240 0.480 1.100 0.660 ;
        RECT  0.920 0.940 1.340 1.220 ;
        RECT  0.920 0.480 1.100 1.480 ;
        RECT  0.100 1.320 1.100 1.480 ;
        RECT  0.100 1.320 0.380 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END ND4B1M0HM

MACRO ND3M8HM
    CLASS CORE ;
    FOREIGN ND3M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.442  LAYER ME1  ;
        ANTENNAGATEAREA 0.442  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.554  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.120 2.700 1.320 ;
        LAYER ME2 ;
        RECT  2.440 0.840 2.760 1.380 ;
        LAYER ME1 ;
        RECT  2.340 1.060 3.340 1.380 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.479  LAYER ME1  ;
        ANTENNAGATEAREA 0.479  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.434  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.120 4.300 1.320 ;
        LAYER ME2 ;
        RECT  4.040 0.840 4.360 1.380 ;
        LAYER ME1 ;
        RECT  3.900 1.060 4.900 1.380 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.442  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.060 1.820 1.380 ;
        RECT  0.440 0.840 0.700 1.380 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.637  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.540 5.500 1.740 ;
        RECT  5.240 0.660 5.500 1.740 ;
        RECT  3.980 0.660 5.500 0.820 ;
        RECT  4.580 1.540 4.780 1.960 ;
        RECT  3.540 1.540 3.740 1.960 ;
        RECT  2.500 1.540 2.700 1.960 ;
        RECT  1.460 1.540 1.660 1.960 ;
        RECT  0.420 1.540 0.620 1.960 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.060 1.900 5.340 2.540 ;
        RECT  4.020 1.900 4.300 2.540 ;
        RECT  2.980 1.900 3.260 2.540 ;
        RECT  1.940 1.900 2.220 2.540 ;
        RECT  0.900 1.900 1.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  1.420 -0.140 1.700 0.500 ;
        RECT  0.420 -0.140 0.620 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.900 0.370 1.120 0.820 ;
        RECT  0.900 0.660 3.300 0.820 ;
        RECT  2.460 0.300 5.900 0.500 ;
        RECT  5.680 0.300 5.900 0.580 ;
        LAYER VTPH ;
        RECT  5.570 1.140 6.000 2.400 ;
        RECT  0.000 1.230 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
        RECT  0.000 0.000 5.570 1.230 ;
    END
END ND3M8HM

MACRO ND3M6HM
    CLASS CORE ;
    FOREIGN ND3M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.359  LAYER ME1  ;
        ANTENNAGATEAREA 0.359  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.913  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.120 2.700 1.320 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.500 ;
        LAYER ME1 ;
        RECT  2.060 1.060 3.060 1.380 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.359  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.060 4.620 1.380 ;
        RECT  3.300 0.840 3.500 1.380 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.359  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 1.540 1.380 ;
        RECT  0.100 0.840 0.300 1.380 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.224  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.140 1.540 5.100 1.740 ;
        RECT  4.900 0.360 5.100 1.740 ;
        RECT  3.680 0.660 5.100 0.860 ;
        RECT  4.780 0.360 5.100 0.860 ;
        RECT  4.300 1.540 4.500 2.030 ;
        RECT  3.260 1.540 3.460 2.030 ;
        RECT  2.220 1.540 2.420 2.030 ;
        RECT  1.180 1.540 1.380 2.030 ;
        RECT  0.140 1.540 0.340 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.100 -0.140 0.380 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.390 0.900 0.860 ;
        RECT  1.660 0.360 1.940 0.860 ;
        RECT  0.620 0.660 3.040 0.860 ;
        RECT  2.180 0.300 4.540 0.460 ;
        RECT  2.180 0.300 2.460 0.500 ;
        RECT  4.260 0.300 4.540 0.500 ;
        RECT  3.220 0.300 3.500 0.560 ;
        LAYER VTPH ;
        RECT  0.000 1.380 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.380 ;
    END
END ND3M6HM

MACRO ND3M4HM
    CLASS CORE ;
    FOREIGN ND3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.239  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.080 2.200 1.280 ;
        RECT  1.300 0.840 1.500 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.239  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.670 0.760 3.100 1.280 ;
        RECT  1.660 0.760 3.100 0.920 ;
        RECT  1.660 0.390 1.860 0.920 ;
        RECT  0.800 0.390 1.860 0.590 ;
        RECT  0.800 0.390 1.080 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.239  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.440 3.460 1.600 ;
        RECT  3.260 1.060 3.460 1.600 ;
        RECT  0.100 1.060 0.560 1.600 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.903  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.580 1.760 3.900 1.920 ;
        RECT  3.700 0.680 3.900 1.920 ;
        RECT  3.260 0.680 3.900 0.840 ;
        RECT  3.260 0.340 3.420 0.840 ;
        RECT  2.020 0.340 3.420 0.500 ;
        RECT  2.020 0.340 2.300 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.420 2.080 3.700 2.540 ;
        RECT  2.300 2.080 2.580 2.540 ;
        RECT  1.180 2.080 1.460 2.540 ;
        RECT  0.140 1.760 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.620 -0.140 3.900 0.500 ;
        RECT  0.140 -0.140 0.340 0.670 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END ND3M4HM

MACRO ND3M3HM
    CLASS CORE ;
    FOREIGN ND3M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER ME1  ;
        ANTENNAGATEAREA 0.181  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.411  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.060 1.500 1.260 ;
        LAYER ME2 ;
        RECT  1.300 0.900 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.200 1.050 1.810 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.700 2.320 1.280 ;
        RECT  0.760 0.700 2.320 0.860 ;
        RECT  0.760 0.700 1.040 1.080 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.440 2.740 1.600 ;
        RECT  2.520 1.060 2.740 1.600 ;
        RECT  0.100 0.820 0.500 1.600 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.738  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 1.760 3.100 1.980 ;
        RECT  2.900 0.540 3.100 1.980 ;
        RECT  2.520 0.540 3.100 0.700 ;
        RECT  0.580 1.760 3.100 1.920 ;
        RECT  2.520 0.340 2.680 0.700 ;
        RECT  1.380 0.340 2.680 0.500 ;
        RECT  1.700 1.760 1.980 2.060 ;
        RECT  0.580 1.760 0.860 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.840 -0.140 3.060 0.380 ;
        RECT  0.100 -0.140 0.380 0.500 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END ND3M3HM

MACRO ND3M2HM
    CLASS CORE ;
    FOREIGN ND3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.760 1.640 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.770 1.100 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.680 1.280 ;
        RECT  0.100 1.000 0.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.538  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.540 2.300 1.740 ;
        RECT  2.100 0.300 2.300 1.740 ;
        RECT  1.580 0.300 2.300 0.500 ;
        RECT  1.700 1.540 1.900 2.030 ;
        RECT  0.660 1.540 0.860 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.760 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.260 -0.140 0.460 0.670 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END ND3M2HM

MACRO ND3M1HM
    CLASS CORE ;
    FOREIGN ND3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.640 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.790 1.100 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.680 1.280 ;
        RECT  0.100 1.000 0.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.378  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.540 2.300 1.740 ;
        RECT  2.100 0.480 2.300 1.740 ;
        RECT  1.580 0.480 2.300 0.680 ;
        RECT  1.700 1.540 1.900 2.090 ;
        RECT  0.660 1.540 0.860 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.260 -0.140 0.460 0.710 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END ND3M1HM

MACRO ND3M16HM
    CLASS CORE ;
    FOREIGN ND3M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.946  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 1.140 10.140 1.420 ;
        RECT  7.300 0.840 7.560 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.958  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 1.140 6.760 1.560 ;
        RECT  4.220 1.140 6.760 1.390 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.958  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.140 3.290 1.390 ;
        RECT  0.440 1.140 0.760 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.047  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.300 1.580 10.700 1.900 ;
        RECT  10.500 0.660 10.700 1.900 ;
        RECT  7.860 0.660 10.700 0.820 ;
        RECT  7.260 1.580 10.700 1.740 ;
        RECT  9.340 1.580 9.620 1.890 ;
        RECT  8.300 1.580 8.580 1.890 ;
        RECT  6.100 1.760 7.540 1.920 ;
        RECT  7.260 1.580 7.540 1.920 ;
        RECT  6.100 1.580 6.300 1.920 ;
        RECT  0.940 1.580 6.300 1.740 ;
        RECT  5.100 1.580 5.380 1.870 ;
        RECT  4.060 1.580 4.340 1.870 ;
        RECT  3.020 1.580 3.300 1.870 ;
        RECT  1.980 1.580 2.260 1.870 ;
        RECT  0.940 1.580 1.220 1.870 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  9.860 1.900 10.140 2.540 ;
        RECT  8.820 1.900 9.100 2.540 ;
        RECT  7.780 1.900 8.060 2.540 ;
        RECT  6.700 2.080 6.980 2.540 ;
        RECT  5.620 1.900 5.900 2.540 ;
        RECT  4.580 1.900 4.860 2.540 ;
        RECT  3.540 1.900 3.820 2.540 ;
        RECT  2.500 1.900 2.780 2.540 ;
        RECT  1.460 1.900 1.740 2.540 ;
        RECT  0.420 1.900 0.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.100 -0.140 0.380 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.480 0.860 0.820 ;
        RECT  0.660 0.660 7.140 0.820 ;
        RECT  6.860 0.660 7.140 0.880 ;
        RECT  4.200 0.340 10.840 0.500 ;
        LAYER VTPH ;
        RECT  2.490 1.230 5.030 2.400 ;
        RECT  0.000 1.240 7.100 2.400 ;
        RECT  0.000 1.320 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.230 ;
        RECT  0.000 0.000 2.490 1.240 ;
        RECT  5.030 0.000 11.200 1.240 ;
        RECT  7.100 0.000 11.200 1.320 ;
    END
END ND3M16HM

MACRO ND3M12HM
    CLASS CORE ;
    FOREIGN ND3M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.718  LAYER ME1  ;
        ANTENNAGATEAREA 0.718  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.500 1.150 6.700 1.350 ;
        LAYER ME2 ;
        RECT  6.500 0.840 6.700 1.560 ;
        LAYER ME1 ;
        RECT  5.700 1.140 7.780 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.718  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.100 1.140 5.500 1.360 ;
        RECT  5.240 0.840 5.500 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.718  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.140 2.580 1.360 ;
        RECT  0.500 0.840 0.700 1.360 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.390  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.580 8.300 1.740 ;
        RECT  8.100 0.440 8.300 1.740 ;
        RECT  5.820 0.770 8.300 0.980 ;
        RECT  7.900 0.440 8.300 0.980 ;
        RECT  7.380 1.580 7.660 1.990 ;
        RECT  6.340 1.580 6.620 1.990 ;
        RECT  5.300 1.580 5.580 1.990 ;
        RECT  4.260 1.580 4.540 1.990 ;
        RECT  3.220 1.580 3.500 1.990 ;
        RECT  2.180 1.580 2.460 1.990 ;
        RECT  1.140 1.580 1.420 1.990 ;
        RECT  0.100 1.580 0.380 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.200 -0.140 1.420 0.560 ;
        RECT  0.100 -0.140 0.380 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.370 1.040 0.650 ;
        RECT  2.700 0.520 2.980 0.980 ;
        RECT  0.880 0.370 1.040 0.980 ;
        RECT  1.660 0.520 1.940 0.980 ;
        RECT  2.700 0.760 5.060 0.980 ;
        RECT  0.880 0.780 5.060 0.980 ;
        RECT  3.220 0.370 7.660 0.590 ;
        LAYER VTPH ;
        RECT  8.000 1.140 8.400 2.400 ;
        RECT  0.000 1.290 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
        RECT  0.000 0.000 8.000 1.290 ;
    END
END ND3M12HM

MACRO ND3M0HM
    CLASS CORE ;
    FOREIGN ND3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.066  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.520 0.840 1.900 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.066  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.790 1.160 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.066  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.600 1.280 ;
        RECT  0.100 1.000 0.360 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.347  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 1.500 2.300 2.090 ;
        RECT  2.100 0.460 2.300 2.090 ;
        RECT  1.900 0.460 2.300 0.680 ;
        RECT  0.700 1.500 2.300 1.700 ;
        RECT  0.700 1.500 0.980 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.300 1.860 1.580 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.140 -0.140 0.340 0.750 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END ND3M0HM

MACRO ND3B1M8HM
    CLASS CORE ;
    FOREIGN ND3B1M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.040 1.080 4.360 1.500 ;
        RECT  3.080 1.080 4.360 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.479  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.640 1.080 5.640 1.360 ;
        RECT  4.640 1.080 5.100 1.560 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.240 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.665  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.320 1.540 6.600 1.960 ;
        RECT  5.280 1.540 6.600 1.700 ;
        RECT  6.060 0.700 6.300 1.700 ;
        RECT  4.700 0.700 6.300 0.860 ;
        RECT  3.680 1.720 5.600 1.880 ;
        RECT  5.280 1.540 5.600 1.880 ;
        RECT  3.680 1.540 3.870 1.880 ;
        RECT  1.640 1.540 3.870 1.700 ;
        RECT  2.680 1.540 2.960 1.810 ;
        RECT  1.640 1.540 1.930 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.800 1.900 6.080 2.540 ;
        RECT  4.320 2.080 4.960 2.540 ;
        RECT  3.200 1.900 3.480 2.540 ;
        RECT  2.160 1.900 2.440 2.540 ;
        RECT  1.180 1.690 1.400 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  2.160 -0.140 2.440 0.500 ;
        RECT  1.120 -0.140 1.400 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.410 0.950 0.630 ;
        RECT  0.750 1.120 2.560 1.320 ;
        RECT  0.750 0.410 0.950 1.680 ;
        RECT  0.100 1.480 0.950 1.680 ;
        RECT  0.100 1.480 0.380 2.060 ;
        RECT  1.640 0.470 1.920 0.860 ;
        RECT  1.640 0.660 4.000 0.860 ;
        RECT  3.140 0.340 6.680 0.500 ;
        RECT  6.400 0.340 6.680 0.560 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.020 2.400 ;
        RECT  0.000 1.230 2.080 2.400 ;
        RECT  3.560 1.230 6.800 2.400 ;
        RECT  0.000 1.240 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
        RECT  1.020 0.000 6.800 1.230 ;
        RECT  2.080 0.000 3.560 1.240 ;
    END
END ND3B1M8HM

MACRO ND3B1M4HM
    CLASS CORE ;
    FOREIGN ND3B1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.239  LAYER ME1  ;
        ANTENNAGATEAREA 0.239  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.003  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.040 2.700 1.240 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.500 ;
        LAYER ME1 ;
        RECT  2.160 1.000 2.800 1.280 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.239  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.120 0.660 3.400 1.280 ;
        RECT  1.620 0.660 3.400 0.820 ;
        RECT  1.620 0.660 1.900 1.280 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.840 1.280 ;
        RECT  0.100 0.840 0.360 1.280 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.881  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 1.760 4.300 1.920 ;
        RECT  4.100 0.620 4.300 1.920 ;
        RECT  3.560 0.620 4.300 0.780 ;
        RECT  3.560 0.340 3.720 0.780 ;
        RECT  2.300 0.340 3.720 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 2.080 4.300 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  1.780 2.080 2.060 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.880 -0.140 4.100 0.380 ;
        RECT  0.900 -0.140 1.180 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 0.370 0.740 0.590 ;
        RECT  0.580 0.370 0.740 0.860 ;
        RECT  0.580 0.660 1.260 0.860 ;
        RECT  1.060 0.660 1.260 1.600 ;
        RECT  3.700 1.020 3.900 1.600 ;
        RECT  0.220 1.440 3.900 1.600 ;
        RECT  0.220 1.440 0.420 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END ND3B1M4HM

MACRO ND3B1M2HM
    CLASS CORE ;
    FOREIGN ND3B1M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.730 1.900 1.300 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.730 2.340 1.300 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 1.020 0.840 1.500 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.538  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.420 1.540 2.700 2.030 ;
        RECT  2.500 0.300 2.700 2.030 ;
        RECT  2.340 0.300 2.700 0.560 ;
        RECT  1.420 1.540 2.700 1.740 ;
        RECT  1.420 1.540 1.660 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.820 2.020 1.100 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.940 -0.140 1.220 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.340 0.500 0.620 0.860 ;
        RECT  0.340 0.660 1.200 0.860 ;
        RECT  1.000 1.020 1.440 1.300 ;
        RECT  1.000 0.660 1.200 1.860 ;
        RECT  0.220 1.660 1.200 1.860 ;
        RECT  0.220 1.660 0.500 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND3B1M2HM

MACRO ND3B1M1HM
    CLASS CORE ;
    FOREIGN ND3B1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.730 1.900 1.250 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.730 2.340 1.250 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 1.020 0.840 1.500 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.378  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.420 1.410 2.700 1.960 ;
        RECT  2.500 0.300 2.700 1.960 ;
        RECT  2.340 0.300 2.700 0.560 ;
        RECT  1.420 1.410 2.700 1.610 ;
        RECT  1.420 1.410 1.660 1.960 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.770 2.180 2.540 ;
        RECT  0.820 2.020 1.100 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.940 -0.140 1.220 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.340 0.500 0.620 0.860 ;
        RECT  0.340 0.660 1.200 0.860 ;
        RECT  1.000 0.960 1.440 1.200 ;
        RECT  1.000 0.660 1.200 1.860 ;
        RECT  0.220 1.660 1.200 1.860 ;
        RECT  0.220 1.660 0.500 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND3B1M1HM

MACRO ND3B1M0HM
    CLASS CORE ;
    FOREIGN ND3B1M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.066  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.740 1.920 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.066  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.740 2.340 1.280 ;
        END
    END C
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 1.060 0.840 1.500 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.347  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.360 1.450 2.700 1.730 ;
        RECT  2.500 0.300 2.700 1.730 ;
        RECT  2.340 0.300 2.700 0.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.820 2.030 2.100 2.540 ;
        RECT  0.700 2.030 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  0.940 -0.140 1.220 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.340 0.310 0.620 0.860 ;
        RECT  0.340 0.660 1.200 0.860 ;
        RECT  1.000 0.920 1.360 1.200 ;
        RECT  1.000 0.660 1.200 1.860 ;
        RECT  0.120 1.660 1.200 1.860 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND3B1M0HM

MACRO ND2M8HM
    CLASS CORE ;
    FOREIGN ND2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.502  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 1.150 3.520 1.370 ;
        RECT  0.760 1.440 3.160 1.600 ;
        RECT  2.880 1.150 3.160 1.600 ;
        RECT  0.760 1.150 1.400 1.600 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.502  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.830 3.940 1.300 ;
        RECT  0.280 0.830 3.940 0.990 ;
        RECT  1.880 0.830 2.600 1.270 ;
        RECT  0.280 0.830 0.560 1.300 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.353  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.380 1.540 4.300 1.740 ;
        RECT  4.100 0.510 4.300 1.740 ;
        RECT  0.900 0.510 4.300 0.670 ;
        RECT  0.900 1.760 3.660 1.920 ;
        RECT  3.380 1.540 3.660 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.700 2.080 2.980 2.540 ;
        RECT  1.500 2.080 1.780 2.540 ;
        RECT  0.320 1.540 0.600 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.940 -0.140 4.220 0.350 ;
        RECT  2.100 -0.140 2.380 0.350 ;
        RECT  0.100 -0.140 0.380 0.620 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END ND2M8HM

MACRO ND2M6HM
    CLASS CORE ;
    FOREIGN ND2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.377  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 0.800 2.500 1.100 ;
        RECT  0.100 0.800 2.500 0.960 ;
        RECT  0.100 0.800 0.500 1.350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.377  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.260 3.120 1.420 ;
        RECT  2.840 0.840 3.120 1.420 ;
        RECT  0.760 1.120 1.400 1.420 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.028  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.580 3.500 1.740 ;
        RECT  3.300 0.480 3.500 1.740 ;
        RECT  0.100 0.480 3.500 0.640 ;
        RECT  2.740 1.580 2.940 2.010 ;
        RECT  1.700 1.580 1.900 2.010 ;
        RECT  0.660 1.580 0.860 2.010 ;
        RECT  0.100 0.420 0.380 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.730 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.710 2.400 ;
        RECT  2.680 1.140 3.600 2.400 ;
        RECT  0.000 1.330 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
        RECT  0.710 0.000 2.680 1.330 ;
    END
END ND2M6HM

MACRO ND2M5HM
    CLASS CORE ;
    FOREIGN ND2M5HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.316  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.800 2.320 1.100 ;
        RECT  0.100 0.800 2.320 0.960 ;
        RECT  0.100 0.800 0.500 1.350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.316  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.260 2.740 1.420 ;
        RECT  2.500 0.840 2.740 1.420 ;
        RECT  0.760 1.120 1.400 1.420 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.836  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 1.580 3.100 1.740 ;
        RECT  2.900 0.480 3.100 1.740 ;
        RECT  0.100 0.480 3.100 0.640 ;
        RECT  2.340 1.580 2.540 2.010 ;
        RECT  1.300 1.580 1.500 2.010 ;
        RECT  0.100 0.420 0.380 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 1.900 3.100 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.740 1.900 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.740 -0.140 3.020 0.320 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END ND2M5HM

MACRO ND2M4HM
    CLASS CORE ;
    FOREIGN ND2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.251  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.060 1.500 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.251  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.110 2.280 1.310 ;
        RECT  1.660 0.660 1.860 1.310 ;
        RECT  0.500 0.660 1.860 0.860 ;
        RECT  0.280 1.110 0.700 1.310 ;
        RECT  0.500 0.660 0.700 1.310 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.836  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 1.580 2.700 1.740 ;
        RECT  2.500 0.740 2.700 1.740 ;
        RECT  2.020 0.740 2.700 0.900 ;
        RECT  2.020 0.340 2.180 0.900 ;
        RECT  0.580 1.760 2.020 1.920 ;
        RECT  1.780 1.580 2.020 1.920 ;
        RECT  0.900 0.340 2.180 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        RECT  1.180 2.080 1.460 2.540 ;
        RECT  0.140 1.730 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.340 -0.140 2.540 0.580 ;
        RECT  0.140 -0.140 0.340 0.670 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END ND2M4HM

MACRO ND2M3HM
    CLASS CORE ;
    FOREIGN ND2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.184  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.800 1.400 1.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.184  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.300 1.880 1.500 ;
        RECT  1.600 0.960 1.880 1.500 ;
        RECT  0.280 0.960 0.560 1.500 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.680 2.300 1.880 ;
        RECT  2.100 0.560 2.300 1.880 ;
        RECT  1.560 0.560 2.300 0.760 ;
        RECT  0.940 0.400 1.760 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.820 2.040 2.100 2.540 ;
        RECT  0.740 1.680 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.920 -0.140 2.120 0.400 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.500 1.120 2.400 2.400 ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.120 ;
        RECT  0.000 0.000 0.500 1.140 ;
    END
END ND2M3HM

MACRO ND2M2HM
    CLASS CORE ;
    FOREIGN ND2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.840 1.100 1.380 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.300 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.409  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.700 1.540 1.500 1.740 ;
        RECT  1.300 0.400 1.500 1.740 ;
        RECT  1.020 0.400 1.500 0.680 ;
        RECT  0.700 1.540 0.900 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.180 1.730 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.180 -0.140 0.380 0.670 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END ND2M2HM

MACRO ND2M1HM
    CLASS CORE ;
    FOREIGN ND2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.088  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.840 1.100 1.380 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.088  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.300 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.284  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.700 1.540 1.500 1.740 ;
        RECT  1.300 0.400 1.500 1.740 ;
        RECT  1.020 0.400 1.500 0.680 ;
        RECT  0.700 1.540 0.900 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.180 1.810 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.180 -0.140 0.380 0.680 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END ND2M1HM

MACRO ND2M16HM
    CLASS CORE ;
    FOREIGN ND2M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.998  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.360 6.520 1.520 ;
        RECT  6.240 1.120 6.520 1.520 ;
        RECT  4.280 1.150 4.920 1.520 ;
        RECT  2.520 1.160 3.160 1.520 ;
        RECT  0.760 1.120 1.160 1.520 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.998  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.840 0.800 7.140 1.220 ;
        RECT  0.280 0.800 7.140 0.960 ;
        RECT  5.160 0.800 5.880 1.160 ;
        RECT  3.760 0.800 4.040 1.160 ;
        RECT  1.680 0.800 1.960 1.160 ;
        RECT  0.280 0.800 0.560 1.260 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.509  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 0.480 7.500 1.740 ;
        RECT  6.700 1.580 7.500 1.740 ;
        RECT  0.900 0.480 7.500 0.640 ;
        RECT  0.940 1.720 6.980 1.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  7.220 1.900 7.500 2.540 ;
        RECT  6.140 2.080 6.420 2.540 ;
        RECT  5.020 2.080 5.300 2.540 ;
        RECT  3.880 2.080 4.160 2.540 ;
        RECT  2.660 2.080 2.940 2.540 ;
        RECT  1.540 2.080 1.820 2.540 ;
        RECT  0.420 1.720 0.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.140 -0.140 7.420 0.320 ;
        RECT  5.380 -0.140 5.660 0.320 ;
        RECT  3.580 -0.140 3.860 0.320 ;
        RECT  1.820 -0.140 2.100 0.320 ;
        RECT  0.100 -0.140 0.380 0.620 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END ND2M16HM

MACRO ND2M12HM
    CLASS CORE ;
    FOREIGN ND2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.752  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.800 1.140 5.080 1.420 ;
        RECT  2.440 1.260 5.080 1.420 ;
        RECT  2.440 1.140 3.260 1.420 ;
        RECT  0.860 1.420 2.760 1.590 ;
        RECT  0.860 1.200 1.500 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.752  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.320 0.800 5.540 1.300 ;
        RECT  0.100 0.800 5.540 0.960 ;
        RECT  3.880 0.800 4.180 1.100 ;
        RECT  1.880 0.800 2.160 1.240 ;
        RECT  0.100 0.800 0.500 1.300 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.923  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.020 1.580 5.900 1.740 ;
        RECT  5.700 0.480 5.900 1.740 ;
        RECT  1.000 0.480 5.900 0.640 ;
        RECT  5.090 1.580 5.390 1.900 ;
        RECT  4.040 1.580 4.360 1.900 ;
        RECT  0.580 1.760 3.300 1.920 ;
        RECT  3.020 1.580 3.300 1.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.620 1.900 5.900 2.540 ;
        RECT  4.580 1.900 4.860 2.540 ;
        RECT  3.540 1.900 3.820 2.540 ;
        RECT  2.440 2.080 2.720 2.540 ;
        RECT  1.180 2.080 1.460 2.540 ;
        RECT  0.140 1.680 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.540 -0.140 5.820 0.320 ;
        RECT  3.680 -0.140 3.960 0.320 ;
        RECT  1.920 -0.140 2.200 0.320 ;
        RECT  0.140 -0.140 0.340 0.620 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.730 2.400 ;
        RECT  0.000 1.200 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
        RECT  0.730 0.000 6.000 1.200 ;
    END
END ND2M12HM

MACRO ND2M0HM
    CLASS CORE ;
    FOREIGN ND2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.840 1.100 1.380 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.300 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.540 1.500 1.740 ;
        RECT  1.300 0.400 1.500 1.740 ;
        RECT  1.020 0.400 1.500 0.680 ;
        RECT  0.660 1.540 0.940 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.180 1.840 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.180 -0.140 0.380 0.680 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END ND2M0HM

MACRO ND2B1M8HM
    CLASS CORE ;
    FOREIGN ND2B1M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.502  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.360 1.340 3.960 1.500 ;
        RECT  3.320 1.140 3.960 1.500 ;
        RECT  1.360 1.140 2.000 1.500 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.300 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.224  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 1.700 4.700 1.900 ;
        RECT  4.540 0.500 4.700 1.900 ;
        RECT  1.500 0.500 4.700 0.660 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.380 -0.140 4.660 0.320 ;
        RECT  2.420 -0.140 2.700 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.060 2.080 4.340 2.540 ;
        RECT  2.940 2.080 3.220 2.540 ;
        RECT  1.780 2.080 2.060 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.060 0.680 ;
        RECT  0.860 0.820 4.380 0.980 ;
        RECT  2.200 0.820 2.840 1.180 ;
        RECT  4.160 0.820 4.380 1.220 ;
        RECT  0.860 0.480 1.060 1.710 ;
        RECT  0.100 1.490 1.060 1.710 ;
        RECT  0.100 1.490 0.380 2.090 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END ND2B1M8HM

MACRO ND2B1M4HM
    CLASS CORE ;
    FOREIGN ND2B1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.251  LAYER ME1  ;
        ANTENNAGATEAREA 0.251  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.576  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.120 1.900 1.320 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.560 1.060 2.000 1.380 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.280 1.060 0.760 1.500 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.612  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 1.540 3.100 1.740 ;
        RECT  2.900 0.720 3.100 1.740 ;
        RECT  2.480 0.720 3.100 0.880 ;
        RECT  2.480 0.340 2.640 0.880 ;
        RECT  2.300 1.540 2.500 2.010 ;
        RECT  1.700 0.340 2.640 0.500 ;
        RECT  1.260 1.540 1.460 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.780 1.900 3.060 2.540 ;
        RECT  1.740 1.900 2.020 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.800 -0.140 3.020 0.560 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.310 0.380 0.820 ;
        RECT  0.160 0.660 2.320 0.820 ;
        RECT  2.160 0.660 2.320 1.380 ;
        RECT  2.160 1.100 2.720 1.380 ;
        RECT  0.940 0.660 1.100 1.880 ;
        RECT  0.160 1.720 1.100 1.880 ;
        RECT  0.160 1.720 0.380 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END ND2B1M4HM

MACRO ND2B1M2HM
    CLASS CORE ;
    FOREIGN ND2B1M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.800 1.500 1.380 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.280 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.381  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 1.560 1.900 1.840 ;
        RECT  1.700 0.340 1.900 1.840 ;
        RECT  1.500 0.340 1.900 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.620 1.940 0.820 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.580 -0.140 0.860 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.020 0.680 ;
        RECT  0.860 0.480 1.020 1.680 ;
        RECT  0.100 1.460 1.020 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END ND2B1M2HM

MACRO ND2B1M1HM
    CLASS CORE ;
    FOREIGN ND2B1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.088  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.240 0.800 1.540 1.280 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.280 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.269  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 1.440 1.900 1.720 ;
        RECT  1.700 0.340 1.900 1.720 ;
        RECT  1.500 0.340 1.900 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.580 1.940 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.580 -0.140 0.860 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.020 0.680 ;
        RECT  0.860 0.480 1.020 1.680 ;
        RECT  0.100 1.460 1.020 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END ND2B1M1HM

MACRO ND2B1M12HM
    CLASS CORE ;
    FOREIGN ND2B1M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.752  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 1.380 6.200 1.540 ;
        RECT  5.560 1.120 6.200 1.540 ;
        RECT  3.720 1.120 4.360 1.540 ;
        RECT  1.840 1.120 2.120 1.540 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.251  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 1.080 1.300 ;
        RECT  0.100 0.840 0.360 1.300 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.836  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.700 6.960 1.900 ;
        RECT  6.800 0.480 6.960 1.900 ;
        RECT  1.940 0.480 6.960 0.640 ;
        RECT  1.700 1.700 1.900 2.050 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.700 2.080 6.980 2.540 ;
        RECT  5.580 2.080 5.860 2.540 ;
        RECT  4.460 2.080 4.740 2.540 ;
        RECT  3.340 2.080 3.620 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.690 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.620 -0.140 6.900 0.320 ;
        RECT  4.860 -0.140 5.140 0.320 ;
        RECT  2.940 -0.140 3.220 0.320 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.390 0.860 0.860 ;
        RECT  0.660 0.660 1.560 0.860 ;
        RECT  1.380 0.800 6.640 0.960 ;
        RECT  4.680 0.800 4.960 1.160 ;
        RECT  2.720 0.800 3.360 1.180 ;
        RECT  6.440 0.800 6.640 1.300 ;
        RECT  1.380 0.660 1.540 1.740 ;
        RECT  0.660 1.540 1.540 1.740 ;
        RECT  0.660 1.540 0.860 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END ND2B1M12HM

MACRO ND2B1M0HM
    CLASS CORE ;
    FOREIGN ND2B1M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.240 0.800 1.540 1.280 ;
        END
    END B
    PIN NA
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.044  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.280 ;
        END
    END NA
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.217  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 1.440 1.900 1.720 ;
        RECT  1.700 0.330 1.900 1.720 ;
        RECT  1.500 0.330 1.900 0.590 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.580 1.940 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.580 -0.140 0.860 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.020 0.680 ;
        RECT  0.860 0.480 1.020 1.680 ;
        RECT  0.100 1.460 1.020 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END ND2B1M0HM

MACRO MXB4M4HM
    CLASS CORE ;
    FOREIGN MXB4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.407  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.120 3.100 1.320 ;
        LAYER ME2 ;
        RECT  2.900 0.790 3.100 1.440 ;
        LAYER ME1 ;
        RECT  2.480 1.120 3.480 1.320 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.681  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.020 1.000 5.220 1.200 ;
        LAYER ME2 ;
        RECT  4.900 0.670 5.220 1.320 ;
        LAYER ME1 ;
        RECT  4.920 0.980 5.350 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.100 1.040 8.300 1.560 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.320 1.560 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.272  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.248  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 9.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.000 1.700 1.660 2.080 ;
        RECT  1.000 0.730 1.200 2.080 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 0.980 9.910 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.468  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.100 1.680 13.500 1.880 ;
        RECT  13.300 0.370 13.500 1.880 ;
        RECT  13.100 0.370 13.500 0.570 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.660 1.480 13.860 2.540 ;
        RECT  12.620 1.480 12.820 2.540 ;
        RECT  8.390 2.080 8.670 2.540 ;
        RECT  4.570 2.080 4.850 2.540 ;
        RECT  4.130 2.080 4.410 2.540 ;
        RECT  3.080 1.860 3.360 2.540 ;
        RECT  0.140 1.820 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.660 -0.140 13.860 0.710 ;
        RECT  12.580 -0.140 12.860 0.540 ;
        RECT  9.430 -0.140 9.630 0.380 ;
        RECT  8.480 -0.140 8.700 0.560 ;
        RECT  4.610 -0.140 4.890 0.500 ;
        RECT  2.830 -0.140 3.110 0.320 ;
        RECT  0.140 -0.140 0.340 0.710 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.350 0.840 2.050 ;
        RECT  2.070 0.640 2.350 0.960 ;
        RECT  2.070 0.800 3.960 0.960 ;
        RECT  3.680 0.800 3.960 1.380 ;
        RECT  2.140 0.640 2.300 1.760 ;
        RECT  2.140 1.560 2.600 1.760 ;
        RECT  1.710 0.320 2.670 0.480 ;
        RECT  1.710 0.320 1.910 0.600 ;
        RECT  4.010 0.320 4.290 0.640 ;
        RECT  2.510 0.480 4.290 0.640 ;
        RECT  4.120 0.320 4.290 0.820 ;
        RECT  4.120 0.660 5.670 0.820 ;
        RECT  5.510 0.660 5.670 1.280 ;
        RECT  4.120 0.320 4.280 1.600 ;
        RECT  4.120 1.400 4.440 1.600 ;
        RECT  5.090 0.340 6.110 0.500 ;
        RECT  5.830 0.340 6.110 1.440 ;
        RECT  4.440 1.000 4.760 1.200 ;
        RECT  7.070 0.780 7.230 1.250 ;
        RECT  6.270 1.090 7.230 1.250 ;
        RECT  4.600 1.000 4.760 1.600 ;
        RECT  4.600 1.440 5.490 1.600 ;
        RECT  6.270 1.090 6.430 1.760 ;
        RECT  5.330 1.600 6.430 1.760 ;
        RECT  7.710 0.640 7.990 0.860 ;
        RECT  7.710 0.640 7.910 1.740 ;
        RECT  6.310 0.320 8.320 0.480 ;
        RECT  6.310 0.320 7.550 0.520 ;
        RECT  8.160 0.320 8.320 0.880 ;
        RECT  8.160 0.720 8.750 0.880 ;
        RECT  8.590 0.720 8.750 1.350 ;
        RECT  7.390 0.320 7.550 1.760 ;
        RECT  6.590 1.560 7.550 1.760 ;
        RECT  10.110 0.640 10.390 1.760 ;
        RECT  9.790 0.320 10.870 0.480 ;
        RECT  9.790 0.320 9.950 0.720 ;
        RECT  8.910 0.560 9.950 0.720 ;
        RECT  8.910 0.560 9.100 1.600 ;
        RECT  8.910 1.440 9.310 1.600 ;
        RECT  10.590 0.320 10.870 1.760 ;
        RECT  11.630 0.640 11.990 0.860 ;
        RECT  11.630 0.640 11.910 1.760 ;
        RECT  1.100 0.390 1.550 0.550 ;
        RECT  1.390 0.390 1.550 1.450 ;
        RECT  1.390 1.290 1.980 1.450 ;
        RECT  2.760 1.540 3.680 1.700 ;
        RECT  3.520 1.540 3.680 1.920 ;
        RECT  1.820 1.290 1.980 2.080 ;
        RECT  3.520 1.760 5.170 1.920 ;
        RECT  8.070 1.760 8.990 1.920 ;
        RECT  2.760 1.540 2.920 2.080 ;
        RECT  1.820 1.920 2.920 2.080 ;
        RECT  5.010 1.920 8.230 2.080 ;
        RECT  12.150 1.070 12.350 2.080 ;
        RECT  8.830 1.920 12.350 2.080 ;
        RECT  11.110 0.320 12.310 0.480 ;
        RECT  12.150 0.320 12.310 0.910 ;
        RECT  12.150 0.750 13.140 0.910 ;
        RECT  12.980 0.750 13.140 1.300 ;
        RECT  11.110 0.320 11.390 1.760 ;
        LAYER VTPH ;
        RECT  3.040 0.850 4.260 2.400 ;
        RECT  5.540 0.920 6.410 2.400 ;
        RECT  3.040 1.060 6.410 2.400 ;
        RECT  8.580 1.080 9.840 2.400 ;
        RECT  2.160 1.160 9.840 2.400 ;
        RECT  0.000 1.140 1.040 2.400 ;
        RECT  11.590 1.160 14.000 2.400 ;
        RECT  2.160 1.240 14.000 2.400 ;
        RECT  12.100 1.140 14.000 2.400 ;
        RECT  0.000 1.260 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 0.850 ;
        RECT  4.260 0.000 14.000 0.920 ;
        RECT  4.260 0.000 5.540 1.060 ;
        RECT  6.410 0.000 14.000 1.080 ;
        RECT  0.000 0.000 3.040 1.140 ;
        RECT  9.840 0.000 14.000 1.140 ;
        RECT  1.040 0.000 3.040 1.160 ;
        RECT  6.410 0.000 8.580 1.160 ;
        RECT  9.840 0.000 12.100 1.160 ;
        RECT  9.840 0.000 11.590 1.240 ;
        RECT  1.040 0.000 2.160 1.260 ;
    END
END MXB4M4HM

MACRO MXB4M2HM
    CLASS CORE ;
    FOREIGN MXB4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.194  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.120 3.100 1.320 ;
        LAYER ME2 ;
        RECT  2.900 0.790 3.100 1.440 ;
        LAYER ME1 ;
        RECT  2.480 1.120 3.480 1.320 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.727  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.020 1.000 5.220 1.200 ;
        LAYER ME2 ;
        RECT  4.900 0.670 5.220 1.320 ;
        LAYER ME1 ;
        RECT  4.920 0.980 5.350 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.100 1.040 8.300 1.560 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.320 1.560 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.272  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.254  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 8.932  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.000 1.700 1.660 2.080 ;
        RECT  1.000 0.770 1.200 2.080 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.700 0.980 9.910 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.950 1.680 13.500 1.880 ;
        RECT  13.300 0.400 13.500 1.880 ;
        RECT  12.950 0.400 13.500 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.470 1.480 12.670 2.540 ;
        RECT  8.390 2.080 8.670 2.540 ;
        RECT  4.570 2.080 4.850 2.540 ;
        RECT  4.130 2.080 4.410 2.540 ;
        RECT  3.080 1.860 3.360 2.540 ;
        RECT  0.140 1.820 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.470 -0.140 12.670 0.560 ;
        RECT  9.430 -0.140 9.630 0.380 ;
        RECT  8.480 -0.140 8.680 0.560 ;
        RECT  4.610 -0.140 4.890 0.500 ;
        RECT  2.830 -0.140 3.110 0.320 ;
        RECT  0.140 -0.140 0.340 0.710 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.350 0.840 2.050 ;
        RECT  2.070 0.640 2.350 0.960 ;
        RECT  2.070 0.800 3.960 0.960 ;
        RECT  3.680 0.800 3.960 1.380 ;
        RECT  2.140 0.640 2.300 1.760 ;
        RECT  2.140 1.560 2.600 1.760 ;
        RECT  1.710 0.320 2.670 0.480 ;
        RECT  1.710 0.320 1.910 0.600 ;
        RECT  4.010 0.320 4.290 0.640 ;
        RECT  2.510 0.480 4.290 0.640 ;
        RECT  4.120 0.320 4.290 0.820 ;
        RECT  4.120 0.660 5.670 0.820 ;
        RECT  5.510 0.660 5.670 1.280 ;
        RECT  4.120 0.320 4.280 1.600 ;
        RECT  4.120 1.400 4.440 1.600 ;
        RECT  5.090 0.340 6.110 0.500 ;
        RECT  5.830 0.340 6.110 1.440 ;
        RECT  4.440 1.000 4.760 1.200 ;
        RECT  7.070 0.780 7.230 1.250 ;
        RECT  6.270 1.090 7.230 1.250 ;
        RECT  4.600 1.000 4.760 1.600 ;
        RECT  4.600 1.440 5.490 1.600 ;
        RECT  6.270 1.090 6.430 1.760 ;
        RECT  5.330 1.600 6.430 1.760 ;
        RECT  7.710 0.640 7.990 0.860 ;
        RECT  7.710 0.640 7.910 1.740 ;
        RECT  6.310 0.320 8.320 0.480 ;
        RECT  6.310 0.320 7.550 0.520 ;
        RECT  8.160 0.320 8.320 0.880 ;
        RECT  8.160 0.720 8.750 0.880 ;
        RECT  8.590 0.720 8.750 1.350 ;
        RECT  7.390 0.320 7.550 1.760 ;
        RECT  6.590 1.560 7.550 1.760 ;
        RECT  10.110 0.640 10.390 1.760 ;
        RECT  9.790 0.320 10.870 0.480 ;
        RECT  9.790 0.320 9.950 0.720 ;
        RECT  8.910 0.560 9.950 0.720 ;
        RECT  8.910 0.560 9.100 1.600 ;
        RECT  8.910 1.440 9.310 1.600 ;
        RECT  10.590 0.320 10.870 1.760 ;
        RECT  11.630 0.620 11.990 0.840 ;
        RECT  11.630 0.620 11.910 1.760 ;
        RECT  1.100 0.390 1.550 0.550 ;
        RECT  1.390 0.390 1.550 1.450 ;
        RECT  1.390 1.290 1.980 1.450 ;
        RECT  2.760 1.540 3.680 1.700 ;
        RECT  3.520 1.540 3.680 1.920 ;
        RECT  1.820 1.290 1.980 2.080 ;
        RECT  3.520 1.760 5.170 1.920 ;
        RECT  8.070 1.760 8.990 1.920 ;
        RECT  2.760 1.540 2.920 2.080 ;
        RECT  1.820 1.920 2.920 2.080 ;
        RECT  5.010 1.920 8.230 2.080 ;
        RECT  12.090 1.060 12.290 2.080 ;
        RECT  8.830 1.920 12.290 2.080 ;
        RECT  11.110 0.300 12.310 0.460 ;
        RECT  12.150 0.300 12.310 0.900 ;
        RECT  12.150 0.740 12.850 0.900 ;
        RECT  12.650 0.740 12.850 1.250 ;
        RECT  11.110 0.300 11.390 1.760 ;
        LAYER VTPH ;
        RECT  3.040 0.850 4.260 2.400 ;
        RECT  5.540 0.920 6.410 2.400 ;
        RECT  3.040 1.060 6.410 2.400 ;
        RECT  8.580 1.080 9.840 2.400 ;
        RECT  2.160 1.160 9.840 2.400 ;
        RECT  0.000 1.140 1.040 2.400 ;
        RECT  2.160 1.240 13.600 2.400 ;
        RECT  11.610 1.140 13.600 2.400 ;
        RECT  0.000 1.260 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 0.850 ;
        RECT  4.260 0.000 13.600 0.920 ;
        RECT  4.260 0.000 5.540 1.060 ;
        RECT  6.410 0.000 13.600 1.080 ;
        RECT  0.000 0.000 3.040 1.140 ;
        RECT  9.840 0.000 13.600 1.140 ;
        RECT  1.040 0.000 3.040 1.160 ;
        RECT  6.410 0.000 8.580 1.160 ;
        RECT  9.840 0.000 11.610 1.240 ;
        RECT  1.040 0.000 2.160 1.260 ;
    END
END MXB4M2HM

MACRO MXB4M1HM
    CLASS CORE ;
    FOREIGN MXB4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.656  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.330 0.970 4.530 1.170 ;
        LAYER ME2 ;
        RECT  4.330 0.840 4.700 1.350 ;
        LAYER ME1 ;
        RECT  4.230 0.940 4.650 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.376  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.150 1.100 7.350 1.300 ;
        LAYER ME2 ;
        RECT  7.090 0.840 7.500 1.400 ;
        LAYER ME1 ;
        RECT  7.090 1.040 7.450 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.940 1.100 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.840 4.050 1.220 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.839  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.256  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 11.108  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.940 2.030 2.100 ;
        RECT  1.870 1.240 2.030 2.100 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  0.500 1.760 1.300 1.920 ;
        RECT  0.500 1.240 0.700 1.920 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.155  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.500 1.150 10.750 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.341  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.080 0.670 9.360 1.780 ;
        RECT  8.900 1.240 9.360 1.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.720 1.740 10.920 2.540 ;
        RECT  7.510 1.840 7.720 2.540 ;
        RECT  4.030 2.080 4.310 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.720 -0.140 10.920 0.840 ;
        RECT  7.630 -0.140 7.830 0.560 ;
        RECT  4.030 -0.140 4.310 0.320 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.430 0.620 1.710 1.660 ;
        RECT  3.030 0.620 3.310 0.840 ;
        RECT  3.030 0.620 3.210 1.780 ;
        RECT  3.370 1.010 3.530 1.600 ;
        RECT  3.370 1.440 5.150 1.600 ;
        RECT  4.790 0.620 5.850 0.780 ;
        RECT  5.310 0.620 5.850 0.820 ;
        RECT  5.310 0.620 5.510 1.780 ;
        RECT  1.100 0.300 3.630 0.460 ;
        RECT  4.470 0.300 6.210 0.460 ;
        RECT  3.470 0.300 3.630 0.640 ;
        RECT  4.470 0.300 4.630 0.640 ;
        RECT  3.470 0.480 4.630 0.640 ;
        RECT  1.100 0.300 1.260 0.700 ;
        RECT  0.140 0.540 1.260 0.700 ;
        RECT  1.870 0.300 2.030 1.070 ;
        RECT  6.010 0.300 6.210 1.350 ;
        RECT  2.650 0.300 2.850 1.560 ;
        RECT  0.140 0.540 0.340 2.050 ;
        RECT  6.750 0.620 7.150 0.840 ;
        RECT  6.750 0.620 6.910 1.780 ;
        RECT  6.750 1.580 7.030 1.780 ;
        RECT  8.560 0.650 8.840 0.850 ;
        RECT  7.190 1.520 8.040 1.680 ;
        RECT  3.390 1.760 4.630 1.920 ;
        RECT  2.190 0.620 2.470 2.100 ;
        RECT  4.470 1.760 4.630 2.100 ;
        RECT  7.880 1.520 8.040 2.100 ;
        RECT  8.560 0.650 8.720 2.100 ;
        RECT  3.390 1.760 3.550 2.100 ;
        RECT  2.190 1.940 3.550 2.100 ;
        RECT  7.190 1.520 7.350 2.100 ;
        RECT  4.470 1.940 7.350 2.100 ;
        RECT  9.660 1.590 9.820 2.100 ;
        RECT  7.880 1.940 9.820 2.100 ;
        RECT  6.390 0.300 7.470 0.460 ;
        RECT  8.210 0.300 9.820 0.460 ;
        RECT  7.310 0.300 7.470 0.880 ;
        RECT  7.310 0.720 8.400 0.880 ;
        RECT  9.660 0.300 9.820 0.960 ;
        RECT  6.390 0.300 6.590 1.780 ;
        RECT  5.830 1.620 6.590 1.780 ;
        RECT  8.210 0.300 8.400 1.780 ;
        RECT  8.200 0.720 8.400 1.780 ;
        RECT  9.520 1.190 10.320 1.390 ;
        RECT  10.120 0.560 10.320 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.950 2.400 ;
        RECT  6.700 1.140 7.840 2.400 ;
        RECT  0.000 1.200 5.730 2.400 ;
        RECT  6.700 1.200 8.630 2.400 ;
        RECT  10.280 1.140 11.200 2.400 ;
        RECT  0.000 1.260 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
        RECT  4.950 0.000 6.700 1.200 ;
        RECT  7.840 0.000 10.280 1.200 ;
        RECT  5.730 0.000 6.700 1.260 ;
        RECT  8.630 0.000 10.280 1.260 ;
    END
END MXB4M1HM

MACRO MXB4M0HM
    CLASS CORE ;
    FOREIGN MXB4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.921  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.330 0.970 4.530 1.170 ;
        LAYER ME2 ;
        RECT  4.330 0.840 4.700 1.350 ;
        LAYER ME1 ;
        RECT  4.230 0.940 4.650 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.508  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.150 1.100 7.350 1.300 ;
        LAYER ME2 ;
        RECT  7.150 0.840 7.500 1.400 ;
        LAYER ME1 ;
        RECT  7.090 1.040 7.450 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.940 1.100 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.840 4.050 1.220 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.839  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.210  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 13.520  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.940 2.030 2.100 ;
        RECT  1.870 1.240 2.030 2.100 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  0.500 1.760 1.300 1.920 ;
        RECT  0.500 1.240 0.700 1.920 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.133  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.500 1.150 10.750 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.256  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.080 0.670 9.360 1.780 ;
        RECT  8.900 1.240 9.360 1.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.720 1.740 10.920 2.540 ;
        RECT  7.510 1.840 7.720 2.540 ;
        RECT  4.030 2.080 4.310 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.720 -0.140 10.920 0.840 ;
        RECT  7.630 -0.140 7.830 0.560 ;
        RECT  4.030 -0.140 4.310 0.320 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.430 0.620 1.710 1.660 ;
        RECT  3.030 0.620 3.310 0.840 ;
        RECT  3.030 0.620 3.210 1.780 ;
        RECT  3.370 1.010 3.530 1.600 ;
        RECT  3.370 1.440 5.150 1.600 ;
        RECT  4.790 0.620 5.850 0.780 ;
        RECT  5.310 0.620 5.850 0.820 ;
        RECT  5.310 0.620 5.510 1.780 ;
        RECT  1.100 0.300 3.630 0.460 ;
        RECT  4.470 0.300 6.210 0.460 ;
        RECT  3.470 0.300 3.630 0.640 ;
        RECT  4.470 0.300 4.630 0.640 ;
        RECT  3.470 0.480 4.630 0.640 ;
        RECT  1.100 0.300 1.260 0.700 ;
        RECT  0.140 0.540 1.260 0.700 ;
        RECT  1.870 0.300 2.030 1.070 ;
        RECT  6.010 0.300 6.210 1.350 ;
        RECT  2.650 0.300 2.850 1.560 ;
        RECT  0.140 0.540 0.340 2.050 ;
        RECT  6.750 0.620 7.150 0.840 ;
        RECT  6.750 0.620 6.910 1.780 ;
        RECT  6.750 1.580 7.030 1.780 ;
        RECT  8.560 0.650 8.840 0.850 ;
        RECT  7.190 1.520 8.040 1.680 ;
        RECT  3.390 1.760 4.630 1.920 ;
        RECT  2.190 0.620 2.470 2.100 ;
        RECT  4.470 1.760 4.630 2.100 ;
        RECT  7.880 1.520 8.040 2.100 ;
        RECT  8.560 0.650 8.720 2.100 ;
        RECT  3.390 1.760 3.550 2.100 ;
        RECT  2.190 1.940 3.550 2.100 ;
        RECT  7.190 1.520 7.350 2.100 ;
        RECT  4.470 1.940 7.350 2.100 ;
        RECT  9.660 1.590 9.820 2.100 ;
        RECT  7.880 1.940 9.820 2.100 ;
        RECT  6.390 0.300 7.470 0.460 ;
        RECT  8.210 0.300 9.820 0.460 ;
        RECT  7.310 0.300 7.470 0.880 ;
        RECT  7.310 0.720 8.400 0.880 ;
        RECT  9.660 0.300 9.820 0.930 ;
        RECT  6.390 0.300 6.590 1.780 ;
        RECT  5.830 1.620 6.590 1.780 ;
        RECT  8.210 0.300 8.400 1.780 ;
        RECT  8.200 0.720 8.400 1.780 ;
        RECT  9.520 1.190 10.320 1.390 ;
        RECT  10.120 0.560 10.320 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.950 2.400 ;
        RECT  6.700 1.140 7.840 2.400 ;
        RECT  0.000 1.200 5.730 2.400 ;
        RECT  6.700 1.200 8.630 2.400 ;
        RECT  10.280 1.140 11.200 2.400 ;
        RECT  0.000 1.260 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
        RECT  4.950 0.000 6.700 1.200 ;
        RECT  7.840 0.000 10.280 1.200 ;
        RECT  5.730 0.000 6.700 1.260 ;
        RECT  8.630 0.000 10.280 1.260 ;
    END
END MXB4M0HM

MACRO MXB3M4HM
    CLASS CORE ;
    FOREIGN MXB3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.180 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 0.840 3.500 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 0.750 6.700 1.160 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.000 1.920 1.900 2.080 ;
        RECT  1.700 1.190 1.900 2.080 ;
        RECT  1.000 1.700 1.160 2.080 ;
        RECT  0.500 1.700 1.160 1.900 ;
        RECT  0.500 0.920 0.660 1.900 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.840 3.940 1.360 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.468  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.080 0.420 8.360 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.640 1.480 8.840 2.540 ;
        RECT  7.600 1.480 7.800 2.540 ;
        RECT  6.520 2.080 6.800 2.540 ;
        RECT  3.620 1.840 3.820 2.540 ;
        RECT  0.550 2.080 0.830 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.640 -0.140 8.840 0.660 ;
        RECT  7.600 -0.140 7.800 0.660 ;
        RECT  6.520 -0.140 6.720 0.560 ;
        RECT  3.460 -0.140 3.660 0.610 ;
        RECT  0.580 -0.140 0.860 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.640 1.620 0.860 ;
        RECT  1.340 0.640 1.540 1.760 ;
        RECT  1.020 0.320 2.760 0.480 ;
        RECT  0.140 0.480 1.180 0.640 ;
        RECT  1.780 0.320 1.940 1.030 ;
        RECT  2.560 0.320 2.760 1.560 ;
        RECT  0.140 0.480 0.340 1.740 ;
        RECT  2.940 0.390 3.140 1.760 ;
        RECT  4.480 0.640 4.840 0.800 ;
        RECT  3.300 1.520 4.150 1.680 ;
        RECT  4.680 0.640 4.840 2.080 ;
        RECT  2.100 0.640 2.380 2.080 ;
        RECT  3.980 1.520 4.150 2.080 ;
        RECT  3.300 1.520 3.460 2.080 ;
        RECT  2.100 1.920 3.460 2.080 ;
        RECT  4.680 1.800 4.990 2.080 ;
        RECT  3.980 1.920 4.990 2.080 ;
        RECT  4.100 0.320 5.800 0.480 ;
        RECT  4.100 0.320 4.260 1.140 ;
        RECT  4.100 0.960 4.510 1.140 ;
        RECT  5.580 0.320 5.800 1.560 ;
        RECT  4.310 0.960 4.510 1.740 ;
        RECT  5.960 0.440 6.160 1.600 ;
        RECT  5.960 1.380 6.240 1.600 ;
        RECT  5.120 0.640 5.400 0.860 ;
        RECT  6.880 0.900 7.040 1.550 ;
        RECT  6.400 1.390 7.040 1.550 ;
        RECT  5.240 0.640 5.400 1.920 ;
        RECT  6.400 1.390 6.560 1.920 ;
        RECT  5.240 1.760 6.560 1.920 ;
        RECT  7.080 0.420 7.360 0.620 ;
        RECT  7.200 0.980 7.920 1.180 ;
        RECT  7.200 0.420 7.360 1.970 ;
        RECT  7.080 1.770 7.360 1.970 ;
        LAYER VTPH ;
        RECT  5.630 1.080 7.550 2.400 ;
        RECT  0.000 1.140 1.090 2.400 ;
        RECT  5.630 1.140 9.200 2.400 ;
        RECT  0.000 1.160 9.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.200 1.080 ;
        RECT  0.000 0.000 5.630 1.140 ;
        RECT  7.550 0.000 9.200 1.140 ;
        RECT  1.090 0.000 5.630 1.160 ;
    END
END MXB3M4HM

MACRO MXB3M2HM
    CLASS CORE ;
    FOREIGN MXB3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.180 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 0.840 3.500 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 0.750 6.700 1.160 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.000 1.940 1.900 2.100 ;
        RECT  1.700 1.280 1.900 2.100 ;
        RECT  1.000 1.700 1.160 2.100 ;
        RECT  0.500 1.700 1.160 1.900 ;
        RECT  0.500 0.920 0.660 1.900 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.840 3.940 1.360 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.080 0.420 8.360 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.600 1.480 7.800 2.540 ;
        RECT  6.520 2.080 6.800 2.540 ;
        RECT  3.620 1.840 3.820 2.540 ;
        RECT  0.550 2.080 0.830 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.600 -0.140 7.800 0.660 ;
        RECT  6.520 -0.140 6.720 0.560 ;
        RECT  3.460 -0.140 3.660 0.610 ;
        RECT  0.580 -0.140 0.860 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.620 1.620 0.840 ;
        RECT  1.340 0.620 1.540 1.760 ;
        RECT  1.020 0.300 2.760 0.460 ;
        RECT  1.020 0.300 1.180 0.640 ;
        RECT  0.140 0.480 1.180 0.640 ;
        RECT  1.780 0.300 1.940 1.120 ;
        RECT  2.560 0.300 2.760 1.560 ;
        RECT  0.140 0.480 0.340 1.720 ;
        RECT  2.940 0.390 3.140 1.760 ;
        RECT  4.480 0.620 4.840 0.780 ;
        RECT  3.300 1.520 4.150 1.680 ;
        RECT  4.680 0.620 4.840 2.080 ;
        RECT  2.100 0.620 2.380 2.080 ;
        RECT  3.980 1.520 4.150 2.080 ;
        RECT  3.300 1.520 3.460 2.080 ;
        RECT  2.100 1.920 3.460 2.080 ;
        RECT  4.680 1.750 4.990 2.080 ;
        RECT  3.980 1.920 4.990 2.080 ;
        RECT  4.100 0.300 5.800 0.460 ;
        RECT  4.100 0.300 4.260 1.140 ;
        RECT  4.100 0.960 4.510 1.140 ;
        RECT  5.580 0.300 5.800 1.540 ;
        RECT  4.310 0.960 4.510 1.740 ;
        RECT  5.960 0.440 6.160 1.600 ;
        RECT  5.960 1.380 6.240 1.600 ;
        RECT  5.120 0.620 5.400 0.840 ;
        RECT  6.880 0.900 7.040 1.550 ;
        RECT  6.400 1.390 7.040 1.550 ;
        RECT  5.240 0.620 5.400 1.920 ;
        RECT  6.400 1.390 6.560 1.920 ;
        RECT  5.240 1.760 6.560 1.920 ;
        RECT  7.080 0.420 7.360 0.620 ;
        RECT  7.200 0.980 7.920 1.180 ;
        RECT  7.200 0.420 7.360 1.970 ;
        RECT  7.080 1.770 7.360 1.970 ;
        LAYER VTPH ;
        RECT  5.630 1.080 7.400 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.080 ;
        RECT  0.000 0.000 5.630 1.140 ;
        RECT  7.400 0.000 8.800 1.140 ;
    END
END MXB3M2HM

MACRO MXB3M1HM
    CLASS CORE ;
    FOREIGN MXB3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.150 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.270 0.840 3.550 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.790 0.840 7.100 1.250 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.950 1.940 1.910 2.100 ;
        RECT  1.750 1.240 1.910 2.100 ;
        RECT  0.950 1.760 1.110 2.100 ;
        RECT  0.500 1.760 1.110 1.920 ;
        RECT  0.500 0.940 0.700 1.920 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.670 1.080 5.900 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.722  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.300 1.720 5.950 2.000 ;
        RECT  5.350 0.620 5.630 0.840 ;
        RECT  5.300 1.600 5.510 2.000 ;
        RECT  5.350 0.620 5.510 2.000 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.830 1.480 7.030 2.540 ;
        RECT  3.590 1.840 3.790 2.540 ;
        RECT  0.510 2.080 0.790 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.830 -0.140 7.030 0.610 ;
        RECT  3.430 -0.140 3.630 0.680 ;
        RECT  0.590 -0.140 0.790 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.310 0.620 1.590 0.840 ;
        RECT  1.310 0.620 1.510 1.780 ;
        RECT  0.950 0.300 2.730 0.460 ;
        RECT  0.950 0.300 1.110 0.700 ;
        RECT  0.140 0.540 1.110 0.700 ;
        RECT  1.750 0.300 1.910 1.070 ;
        RECT  2.530 0.300 2.730 1.560 ;
        RECT  0.140 0.540 0.340 1.720 ;
        RECT  2.910 0.400 3.110 1.720 ;
        RECT  2.070 0.620 2.350 0.840 ;
        RECT  3.270 1.520 4.110 1.680 ;
        RECT  4.590 0.620 4.870 2.100 ;
        RECT  3.950 1.520 4.110 2.100 ;
        RECT  2.070 0.620 2.230 2.100 ;
        RECT  3.270 1.520 3.430 2.100 ;
        RECT  2.070 1.940 3.430 2.100 ;
        RECT  4.590 1.750 4.930 2.100 ;
        RECT  3.950 1.930 4.930 2.100 ;
        RECT  3.990 0.300 5.950 0.460 ;
        RECT  3.990 0.300 4.430 0.520 ;
        RECT  5.790 0.300 5.950 0.870 ;
        RECT  5.790 0.710 6.310 0.870 ;
        RECT  5.030 0.300 5.190 1.070 ;
        RECT  6.150 0.710 6.310 1.290 ;
        RECT  4.270 0.300 4.430 1.770 ;
        RECT  6.190 0.320 6.630 0.520 ;
        RECT  6.470 0.320 6.630 1.950 ;
        RECT  6.270 1.750 6.630 1.950 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END MXB3M1HM

MACRO MXB3M0HM
    CLASS CORE ;
    FOREIGN MXB3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.150 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.270 0.840 3.550 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.790 0.840 7.100 1.250 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.130  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.990 1.940 1.910 2.100 ;
        RECT  1.750 1.220 1.910 2.100 ;
        RECT  0.990 1.760 1.150 2.100 ;
        RECT  0.500 1.760 1.150 1.920 ;
        RECT  0.500 0.940 0.700 1.920 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.133  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.670 1.080 5.900 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.590  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.300 1.720 5.950 2.000 ;
        RECT  5.350 0.620 5.630 0.840 ;
        RECT  5.300 1.600 5.510 2.000 ;
        RECT  5.350 0.620 5.510 2.000 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.830 1.710 7.030 2.540 ;
        RECT  3.590 1.840 3.790 2.540 ;
        RECT  0.550 2.080 0.830 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.830 -0.140 7.030 0.610 ;
        RECT  3.430 -0.140 3.630 0.680 ;
        RECT  0.590 -0.140 0.790 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.310 0.620 1.590 0.840 ;
        RECT  1.310 0.620 1.510 1.780 ;
        RECT  0.950 0.300 2.730 0.460 ;
        RECT  0.950 0.300 1.110 0.700 ;
        RECT  0.140 0.540 1.110 0.700 ;
        RECT  1.750 0.300 1.910 1.050 ;
        RECT  2.530 0.300 2.730 1.540 ;
        RECT  0.140 0.540 0.340 1.720 ;
        RECT  2.910 0.470 3.110 1.780 ;
        RECT  2.070 0.620 2.350 0.840 ;
        RECT  3.270 1.520 4.110 1.680 ;
        RECT  4.590 0.620 4.870 2.100 ;
        RECT  3.950 1.520 4.110 2.100 ;
        RECT  2.070 0.620 2.230 2.100 ;
        RECT  3.270 1.520 3.430 2.100 ;
        RECT  2.070 1.940 3.430 2.100 ;
        RECT  4.590 1.750 4.930 2.100 ;
        RECT  3.950 1.930 4.930 2.100 ;
        RECT  3.990 0.300 5.950 0.460 ;
        RECT  3.990 0.300 4.430 0.520 ;
        RECT  5.790 0.300 5.950 0.870 ;
        RECT  5.790 0.710 6.310 0.870 ;
        RECT  5.030 0.300 5.190 1.070 ;
        RECT  6.150 0.710 6.310 1.290 ;
        RECT  4.270 0.300 4.430 1.770 ;
        RECT  6.190 0.320 6.630 0.520 ;
        RECT  6.470 0.320 6.630 1.950 ;
        RECT  6.270 1.750 6.630 1.950 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END MXB3M0HM

MACRO MXB2M8HM
    CLASS CORE ;
    FOREIGN MXB2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.145  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.060 1.100 1.260 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.860 0.860 1.200 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.170 1.080 3.510 1.610 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.040 1.940 2.600 2.100 ;
        RECT  2.440 0.760 2.600 2.100 ;
        RECT  1.040 1.660 1.200 2.100 ;
        RECT  0.500 1.660 1.200 1.860 ;
        RECT  0.500 1.020 0.700 1.860 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.090 0.460 6.370 2.100 ;
        RECT  5.150 1.240 6.370 1.560 ;
        RECT  5.050 1.480 5.330 2.100 ;
        RECT  5.150 0.460 5.330 2.100 ;
        RECT  5.050 0.460 5.330 0.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.610 1.480 6.890 2.540 ;
        RECT  5.570 1.850 5.850 2.540 ;
        RECT  4.530 1.520 4.810 2.540 ;
        RECT  3.490 1.880 3.770 2.540 ;
        RECT  0.660 2.020 0.880 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.610 -0.140 6.890 0.740 ;
        RECT  5.570 -0.140 5.850 0.740 ;
        RECT  4.530 -0.140 4.810 0.740 ;
        RECT  3.550 -0.140 3.770 0.590 ;
        RECT  0.660 -0.140 0.880 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.360 0.620 1.640 1.780 ;
        RECT  1.040 0.300 1.960 0.460 ;
        RECT  1.040 0.300 1.200 0.700 ;
        RECT  0.100 0.540 1.200 0.700 ;
        RECT  1.800 0.300 1.960 1.240 ;
        RECT  0.100 0.480 0.330 1.810 ;
        RECT  2.810 0.620 3.010 2.040 ;
        RECT  2.810 1.840 3.170 2.040 ;
        RECT  2.120 0.300 3.350 0.460 ;
        RECT  3.190 0.300 3.350 0.910 ;
        RECT  3.190 0.750 3.830 0.910 ;
        RECT  3.670 0.750 3.830 1.280 ;
        RECT  2.120 0.300 2.280 1.780 ;
        RECT  1.900 1.560 2.280 1.780 ;
        RECT  4.010 1.030 4.970 1.310 ;
        RECT  4.010 0.310 4.290 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.540 2.400 ;
        RECT  3.260 1.140 7.200 2.400 ;
        RECT  0.000 1.200 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
        RECT  2.540 0.000 3.260 1.200 ;
    END
END MXB2M8HM

MACRO MXB2M6HM
    CLASS CORE ;
    FOREIGN MXB2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.145  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.060 1.100 1.260 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.860 0.860 1.200 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.170 1.080 3.510 1.610 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.040 1.940 2.600 2.100 ;
        RECT  2.440 0.760 2.600 2.100 ;
        RECT  1.040 1.660 1.200 2.100 ;
        RECT  0.500 1.660 1.200 1.860 ;
        RECT  0.500 1.020 0.700 1.860 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.090 0.460 6.370 2.100 ;
        RECT  5.150 1.250 6.370 1.560 ;
        RECT  5.050 1.480 5.330 2.100 ;
        RECT  5.150 0.460 5.330 2.100 ;
        RECT  5.050 0.460 5.330 0.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.570 1.850 5.850 2.540 ;
        RECT  4.530 1.820 4.810 2.540 ;
        RECT  3.490 1.880 3.770 2.540 ;
        RECT  0.660 2.020 0.880 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.570 -0.140 5.850 0.740 ;
        RECT  4.530 -0.140 4.810 0.600 ;
        RECT  3.550 -0.140 3.770 0.590 ;
        RECT  0.660 -0.140 0.880 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.360 0.620 1.640 1.780 ;
        RECT  1.040 0.300 1.960 0.460 ;
        RECT  1.040 0.300 1.200 0.700 ;
        RECT  0.100 0.540 1.200 0.700 ;
        RECT  1.800 0.300 1.960 1.240 ;
        RECT  0.100 0.480 0.330 1.810 ;
        RECT  2.810 0.620 3.010 2.040 ;
        RECT  2.810 1.840 3.170 2.040 ;
        RECT  2.120 0.300 3.350 0.460 ;
        RECT  3.190 0.300 3.350 0.910 ;
        RECT  3.190 0.750 3.830 0.910 ;
        RECT  3.670 0.750 3.830 1.280 ;
        RECT  2.120 0.300 2.280 1.780 ;
        RECT  1.900 1.560 2.280 1.780 ;
        RECT  4.010 1.030 4.970 1.310 ;
        RECT  4.010 0.310 4.290 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.540 2.400 ;
        RECT  3.260 1.140 6.800 2.400 ;
        RECT  0.000 1.200 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
        RECT  2.540 0.000 3.260 1.200 ;
    END
END MXB2M6HM

MACRO MXB2M4HM
    CLASS CORE ;
    FOREIGN MXB2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.699  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.060 1.100 1.260 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.860 0.860 1.200 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.170 1.080 3.510 1.610 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.170  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.040 1.940 2.600 2.100 ;
        RECT  2.440 0.760 2.600 2.100 ;
        RECT  1.040 1.660 1.200 2.100 ;
        RECT  0.500 1.660 1.200 1.860 ;
        RECT  0.500 1.020 0.700 1.860 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.150 1.130 5.560 1.560 ;
        RECT  5.050 1.480 5.330 2.100 ;
        RECT  5.150 0.460 5.330 2.100 ;
        RECT  5.050 0.460 5.330 0.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.570 1.850 5.850 2.540 ;
        RECT  4.530 1.820 4.810 2.540 ;
        RECT  3.490 1.880 3.770 2.540 ;
        RECT  0.660 2.020 0.880 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.570 -0.140 5.850 0.740 ;
        RECT  4.530 -0.140 4.810 0.560 ;
        RECT  3.550 -0.140 3.770 0.560 ;
        RECT  0.660 -0.140 0.880 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.360 0.620 1.640 1.780 ;
        RECT  1.040 0.300 1.960 0.460 ;
        RECT  1.040 0.300 1.200 0.700 ;
        RECT  0.100 0.540 1.200 0.700 ;
        RECT  1.800 0.300 1.960 1.240 ;
        RECT  0.100 0.480 0.330 1.810 ;
        RECT  2.810 0.620 3.010 2.040 ;
        RECT  2.810 1.840 3.230 2.040 ;
        RECT  2.120 0.300 3.350 0.460 ;
        RECT  3.190 0.300 3.350 0.910 ;
        RECT  3.190 0.750 3.830 0.910 ;
        RECT  3.670 0.750 3.830 1.280 ;
        RECT  2.120 0.300 2.280 1.780 ;
        RECT  1.900 1.560 2.280 1.780 ;
        RECT  4.010 1.030 4.970 1.310 ;
        RECT  4.010 0.310 4.290 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.540 2.400 ;
        RECT  3.260 1.140 6.000 2.400 ;
        RECT  0.000 1.200 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
        RECT  2.540 0.000 3.260 1.200 ;
    END
END MXB2M4HM

MACRO MXB2M3HM
    CLASS CORE ;
    FOREIGN MXB2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.699  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.060 1.100 1.260 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.860 0.860 1.200 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.170 1.080 3.510 1.610 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.170  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.040 1.940 2.600 2.100 ;
        RECT  2.440 0.760 2.600 2.100 ;
        RECT  1.040 1.660 1.200 2.100 ;
        RECT  0.500 1.660 1.200 1.860 ;
        RECT  0.500 1.020 0.700 1.860 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.376  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.150 0.900 5.560 1.560 ;
        RECT  5.050 1.480 5.330 2.100 ;
        RECT  5.150 0.350 5.330 2.100 ;
        RECT  5.050 0.350 5.330 0.630 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.570 1.850 5.850 2.540 ;
        RECT  4.530 1.820 4.810 2.540 ;
        RECT  3.490 1.880 3.770 2.540 ;
        RECT  0.660 2.020 0.880 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.570 -0.140 5.850 0.630 ;
        RECT  4.530 -0.140 4.810 0.560 ;
        RECT  3.550 -0.140 3.770 0.560 ;
        RECT  0.660 -0.140 0.880 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.360 0.620 1.640 1.780 ;
        RECT  1.040 0.300 1.960 0.460 ;
        RECT  1.040 0.300 1.200 0.700 ;
        RECT  0.100 0.540 1.200 0.700 ;
        RECT  1.800 0.300 1.960 1.240 ;
        RECT  0.100 0.480 0.330 1.810 ;
        RECT  2.810 0.620 3.010 2.040 ;
        RECT  2.810 1.840 3.230 2.040 ;
        RECT  2.120 0.300 3.350 0.460 ;
        RECT  3.190 0.300 3.350 0.910 ;
        RECT  3.190 0.750 3.830 0.910 ;
        RECT  3.670 0.750 3.830 1.280 ;
        RECT  2.120 0.300 2.280 1.780 ;
        RECT  1.900 1.560 2.280 1.780 ;
        RECT  4.010 1.030 4.970 1.310 ;
        RECT  4.010 0.310 4.290 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.540 2.400 ;
        RECT  3.260 1.140 6.000 2.400 ;
        RECT  0.000 1.200 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
        RECT  2.540 0.000 3.260 1.200 ;
    END
END MXB2M3HM

MACRO MXB2M2HM
    CLASS CORE ;
    FOREIGN MXB2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.300 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.880 1.230 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.173  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.060 1.940 2.280 2.100 ;
        RECT  2.120 0.700 2.280 2.100 ;
        RECT  1.060 1.480 1.220 2.100 ;
        RECT  0.500 1.480 1.220 1.640 ;
        RECT  0.500 1.010 0.700 1.640 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.606  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 1.560 1.960 1.720 ;
        RECT  1.780 0.360 1.960 1.720 ;
        RECT  1.640 0.360 1.960 0.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.860 1.610 3.060 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.860 -0.140 3.060 0.610 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.480 1.480 0.680 ;
        RECT  1.320 0.480 1.480 1.180 ;
        RECT  1.320 0.900 1.620 1.180 ;
        RECT  0.140 0.480 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MXB2M2HM

MACRO MXB2M1HM
    CLASS CORE ;
    FOREIGN MXB2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.090  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.800 1.160 1.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.880 1.230 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.060 1.940 2.280 2.100 ;
        RECT  2.120 0.700 2.280 2.100 ;
        RECT  1.060 1.360 1.220 2.100 ;
        RECT  0.500 1.360 1.220 1.520 ;
        RECT  0.500 0.840 0.700 1.520 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.511  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 1.560 1.960 1.720 ;
        RECT  1.780 0.360 1.960 1.720 ;
        RECT  1.640 0.360 1.960 0.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.860 1.610 3.060 2.540 ;
        RECT  0.700 1.680 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.860 -0.140 3.060 0.610 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.480 1.480 0.640 ;
        RECT  1.320 0.480 1.480 1.180 ;
        RECT  1.320 0.900 1.620 1.180 ;
        RECT  0.140 0.360 0.340 1.850 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MXB2M1HM

MACRO MXB2M0HM
    CLASS CORE ;
    FOREIGN MXB2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.840 1.240 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.580 0.800 3.100 1.160 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.980 1.940 2.380 2.100 ;
        RECT  2.160 0.800 2.380 2.100 ;
        RECT  0.980 1.600 1.140 2.100 ;
        RECT  0.490 1.600 1.140 1.760 ;
        RECT  0.490 1.000 0.700 1.760 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.494  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 0.420 2.120 0.640 ;
        RECT  1.540 1.300 2.000 1.780 ;
        RECT  1.840 0.420 2.000 1.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 1.630 3.100 2.540 ;
        RECT  0.390 2.020 0.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.640 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 0.380 0.680 ;
        RECT  0.100 0.500 1.680 0.680 ;
        RECT  1.460 0.500 1.680 1.120 ;
        RECT  0.100 0.340 0.330 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MXB2M0HM

MACRO MUX4M4HM
    CLASS CORE ;
    FOREIGN MUX4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.866  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.010 8.300 1.210 ;
        LAYER ME2 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  8.100 0.860 8.420 1.360 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER ME1  ;
        ANTENNAGATEAREA 0.169  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.582  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.680 1.010 8.880 1.210 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.880 1.560 ;
        LAYER ME1 ;
        RECT  8.580 0.860 8.920 1.360 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.960 0.440 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.120 3.350 1.280 ;
        RECT  2.500 0.900 2.760 1.280 ;
        RECT  2.440 0.900 2.760 1.100 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.400 1.120 4.900 1.560 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.295  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 1.160 7.100 1.440 ;
        RECT  6.100 0.300 6.300 1.440 ;
        RECT  5.120 0.300 6.300 0.460 ;
        RECT  4.360 0.480 5.280 0.640 ;
        RECT  5.120 0.300 5.280 0.640 ;
        RECT  4.360 0.300 4.520 0.640 ;
        RECT  3.600 0.300 4.520 0.460 ;
        RECT  2.920 0.750 3.760 0.950 ;
        RECT  3.600 0.300 3.760 0.950 ;
        RECT  2.920 0.300 3.080 0.950 ;
        RECT  2.460 0.300 3.080 0.730 ;
        RECT  1.020 0.300 3.080 0.460 ;
        RECT  1.020 0.300 1.180 1.580 ;
        END
    END S0
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.260 1.440 12.700 1.600 ;
        RECT  12.500 0.730 12.700 1.600 ;
        RECT  12.260 0.730 12.700 0.890 ;
        RECT  12.260 1.440 12.460 2.080 ;
        RECT  12.260 0.390 12.460 0.890 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.780 1.840 12.980 2.540 ;
        RECT  11.640 1.550 11.840 2.540 ;
        RECT  8.400 1.840 8.600 2.540 ;
        RECT  4.480 2.080 4.760 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.140 1.810 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.780 -0.140 12.980 0.560 ;
        RECT  11.760 -0.140 11.920 0.660 ;
        RECT  8.400 -0.140 8.600 0.380 ;
        RECT  4.680 -0.140 4.960 0.320 ;
        RECT  3.240 -0.140 3.440 0.560 ;
        RECT  0.140 -0.140 0.340 0.700 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 0.840 2.070 ;
        RECT  1.820 0.620 2.300 0.820 ;
        RECT  1.820 0.620 2.020 1.780 ;
        RECT  1.700 1.550 2.020 1.780 ;
        RECT  3.920 0.620 4.200 0.960 ;
        RECT  3.920 0.800 5.280 0.960 ;
        RECT  5.120 0.800 5.280 1.280 ;
        RECT  5.120 1.000 5.600 1.280 ;
        RECT  2.180 1.230 2.340 1.600 ;
        RECT  3.920 0.620 4.080 1.600 ;
        RECT  2.180 1.440 4.080 1.600 ;
        RECT  3.680 1.440 3.960 1.720 ;
        RECT  5.440 0.620 5.920 0.820 ;
        RECT  5.760 0.620 5.920 1.700 ;
        RECT  5.230 1.500 5.920 1.700 ;
        RECT  7.600 0.620 7.880 1.780 ;
        RECT  6.600 0.300 8.240 0.460 ;
        RECT  8.080 0.300 8.240 0.700 ;
        RECT  8.840 0.300 9.360 0.700 ;
        RECT  8.080 0.540 9.360 0.700 ;
        RECT  6.600 0.300 6.760 1.000 ;
        RECT  6.600 0.840 7.420 1.000 ;
        RECT  9.080 0.300 9.360 1.460 ;
        RECT  7.260 0.840 7.420 1.780 ;
        RECT  6.480 1.620 7.420 1.780 ;
        RECT  10.240 0.620 10.800 0.820 ;
        RECT  1.340 0.620 1.620 0.840 ;
        RECT  8.080 1.520 8.920 1.680 ;
        RECT  10.240 0.620 10.400 1.780 ;
        RECT  8.760 1.620 10.400 1.780 ;
        RECT  2.230 1.760 3.520 1.920 ;
        RECT  4.160 1.760 5.080 1.920 ;
        RECT  1.340 0.620 1.540 2.100 ;
        RECT  1.140 1.810 1.540 2.100 ;
        RECT  4.920 1.760 5.080 2.100 ;
        RECT  3.360 1.920 4.320 2.080 ;
        RECT  2.230 1.760 2.390 2.100 ;
        RECT  1.140 1.940 2.390 2.100 ;
        RECT  8.080 1.520 8.240 2.100 ;
        RECT  4.920 1.940 8.240 2.100 ;
        RECT  11.000 0.620 11.280 1.730 ;
        RECT  10.560 1.450 11.280 1.730 ;
        RECT  10.560 1.450 10.720 2.100 ;
        RECT  8.760 1.940 10.720 2.100 ;
        RECT  9.600 0.300 11.600 0.460 ;
        RECT  11.440 0.300 11.600 1.270 ;
        RECT  11.440 1.070 12.340 1.270 ;
        RECT  9.600 0.300 9.880 1.460 ;
        LAYER VTPH ;
        RECT  8.750 0.940 10.180 2.400 ;
        RECT  0.000 1.140 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 0.940 ;
        RECT  0.000 0.000 8.750 1.140 ;
        RECT  10.180 0.000 13.200 1.140 ;
    END
END MUX4M4HM

MACRO MUX4M2HM
    CLASS CORE ;
    FOREIGN MUX4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.281  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.010 8.300 1.210 ;
        LAYER ME2 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  8.100 0.860 8.420 1.360 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.960 0.440 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.120 3.350 1.280 ;
        RECT  2.500 0.900 2.760 1.280 ;
        RECT  2.440 0.900 2.760 1.100 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.400 1.120 4.900 1.560 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.256  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 1.160 7.100 1.440 ;
        RECT  6.100 0.300 6.300 1.440 ;
        RECT  5.120 0.300 6.300 0.460 ;
        RECT  4.360 0.480 5.280 0.640 ;
        RECT  5.120 0.300 5.280 0.640 ;
        RECT  4.360 0.300 4.520 0.640 ;
        RECT  3.600 0.300 4.520 0.460 ;
        RECT  2.920 0.750 3.760 0.950 ;
        RECT  3.600 0.300 3.760 0.950 ;
        RECT  2.920 0.300 3.080 0.950 ;
        RECT  2.460 0.300 3.080 0.730 ;
        RECT  1.020 0.300 3.080 0.460 ;
        RECT  1.020 0.300 1.180 1.580 ;
        END
    END S0
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.220 1.460 12.700 2.080 ;
        RECT  12.500 0.390 12.700 2.080 ;
        RECT  12.220 0.390 12.700 0.720 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.155  LAYER ME1  ;
        ANTENNAGATEAREA 0.155  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.822  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.680 1.010 8.880 1.210 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.880 1.560 ;
        LAYER ME1 ;
        RECT  8.580 0.860 8.920 1.360 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.640 1.550 11.840 2.540 ;
        RECT  8.400 1.840 8.600 2.540 ;
        RECT  4.480 2.080 4.760 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.140 1.810 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.760 -0.140 11.920 0.660 ;
        RECT  8.400 -0.140 8.600 0.380 ;
        RECT  4.680 -0.140 4.960 0.320 ;
        RECT  3.240 -0.140 3.440 0.560 ;
        RECT  0.140 -0.140 0.340 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 0.840 2.070 ;
        RECT  1.820 0.620 2.300 0.820 ;
        RECT  1.820 0.620 2.020 1.780 ;
        RECT  1.700 1.550 2.020 1.780 ;
        RECT  3.920 0.620 4.200 0.960 ;
        RECT  3.920 0.800 5.280 0.960 ;
        RECT  5.120 0.800 5.280 1.280 ;
        RECT  5.120 1.000 5.600 1.280 ;
        RECT  2.180 1.230 2.340 1.600 ;
        RECT  3.920 0.620 4.080 1.600 ;
        RECT  2.180 1.440 4.080 1.600 ;
        RECT  3.680 1.440 3.960 1.720 ;
        RECT  5.440 0.620 5.920 0.820 ;
        RECT  5.760 0.620 5.920 1.760 ;
        RECT  5.240 1.560 5.920 1.760 ;
        RECT  7.600 0.620 7.920 1.780 ;
        RECT  6.600 0.300 8.240 0.460 ;
        RECT  8.080 0.300 8.240 0.700 ;
        RECT  8.840 0.300 9.360 0.700 ;
        RECT  8.080 0.540 9.360 0.700 ;
        RECT  6.600 0.300 6.760 1.000 ;
        RECT  6.600 0.840 7.420 1.000 ;
        RECT  9.080 0.300 9.360 1.460 ;
        RECT  7.260 0.840 7.420 1.780 ;
        RECT  6.340 1.620 7.420 1.780 ;
        RECT  10.240 0.620 10.800 0.820 ;
        RECT  1.340 0.620 1.620 0.840 ;
        RECT  8.080 1.520 8.920 1.680 ;
        RECT  10.240 0.620 10.400 1.780 ;
        RECT  8.760 1.620 10.400 1.780 ;
        RECT  2.230 1.760 3.520 1.920 ;
        RECT  4.160 1.760 5.080 1.920 ;
        RECT  1.340 0.620 1.540 2.100 ;
        RECT  1.140 1.810 1.540 2.100 ;
        RECT  4.920 1.760 5.080 2.100 ;
        RECT  3.360 1.920 4.320 2.080 ;
        RECT  2.230 1.760 2.390 2.100 ;
        RECT  1.140 1.940 2.390 2.100 ;
        RECT  8.080 1.520 8.240 2.100 ;
        RECT  4.920 1.940 8.240 2.100 ;
        RECT  10.560 1.700 11.280 2.100 ;
        RECT  10.960 0.620 11.280 2.100 ;
        RECT  8.760 1.940 11.280 2.100 ;
        RECT  9.600 0.300 11.600 0.460 ;
        RECT  11.440 0.300 11.600 1.230 ;
        RECT  11.440 1.070 12.180 1.230 ;
        RECT  9.600 0.300 9.880 1.460 ;
        LAYER VTPH ;
        RECT  8.750 0.940 10.180 2.400 ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 0.940 ;
        RECT  0.000 0.000 8.750 1.140 ;
        RECT  10.180 0.000 12.800 1.140 ;
    END
END MUX4M2HM

MACRO MUX4M1HM
    CLASS CORE ;
    FOREIGN MUX4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        ANTENNAGATEAREA 0.154  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.844  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.680 1.010 8.880 1.210 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.880 1.560 ;
        LAYER ME1 ;
        RECT  8.580 0.860 8.920 1.360 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.552  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.010 8.300 1.210 ;
        LAYER ME2 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  8.100 0.860 8.420 1.360 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.960 0.440 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.120 3.350 1.280 ;
        RECT  2.500 0.900 2.760 1.280 ;
        RECT  2.440 0.900 2.760 1.100 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.400 1.120 4.900 1.560 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 1.160 7.100 1.440 ;
        RECT  6.100 0.300 6.300 1.440 ;
        RECT  5.120 0.300 6.300 0.460 ;
        RECT  4.360 0.480 5.280 0.640 ;
        RECT  5.120 0.300 5.280 0.640 ;
        RECT  4.360 0.300 4.520 0.640 ;
        RECT  3.600 0.300 4.520 0.460 ;
        RECT  2.920 0.750 3.760 0.950 ;
        RECT  3.600 0.300 3.760 0.950 ;
        RECT  2.920 0.300 3.080 0.950 ;
        RECT  2.460 0.300 3.080 0.730 ;
        RECT  1.020 0.300 3.080 0.460 ;
        RECT  1.020 0.300 1.180 1.580 ;
        END
    END S0
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.200 1.670 12.700 1.920 ;
        RECT  12.480 0.540 12.700 1.920 ;
        RECT  12.200 0.540 12.700 0.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.640 1.550 11.840 2.540 ;
        RECT  8.400 1.840 8.600 2.540 ;
        RECT  4.480 2.080 4.760 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.140 1.810 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.760 -0.140 11.920 0.780 ;
        RECT  8.400 -0.140 8.600 0.380 ;
        RECT  4.680 -0.140 4.960 0.320 ;
        RECT  3.240 -0.140 3.440 0.560 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 0.840 2.070 ;
        RECT  1.820 0.620 2.300 0.820 ;
        RECT  1.820 0.620 2.020 1.780 ;
        RECT  1.700 1.550 2.020 1.780 ;
        RECT  3.920 0.620 4.200 0.960 ;
        RECT  3.920 0.800 5.280 0.960 ;
        RECT  5.120 0.800 5.280 1.280 ;
        RECT  5.120 1.000 5.600 1.280 ;
        RECT  2.180 1.230 2.340 1.600 ;
        RECT  3.920 0.620 4.080 1.600 ;
        RECT  2.180 1.440 4.080 1.600 ;
        RECT  3.680 1.440 3.960 1.720 ;
        RECT  5.440 0.620 5.920 0.820 ;
        RECT  5.760 0.620 5.920 1.760 ;
        RECT  5.240 1.560 5.920 1.760 ;
        RECT  7.600 0.620 7.920 1.780 ;
        RECT  6.540 0.300 8.240 0.460 ;
        RECT  8.080 0.300 8.240 0.700 ;
        RECT  8.840 0.300 9.360 0.700 ;
        RECT  8.080 0.540 9.360 0.700 ;
        RECT  6.540 0.300 6.820 1.000 ;
        RECT  6.540 0.840 7.420 1.000 ;
        RECT  9.080 0.300 9.360 1.460 ;
        RECT  7.260 0.840 7.420 1.780 ;
        RECT  6.340 1.620 7.420 1.780 ;
        RECT  10.240 0.620 10.800 0.820 ;
        RECT  1.340 0.620 1.620 0.840 ;
        RECT  8.080 1.520 8.920 1.680 ;
        RECT  10.240 0.620 10.400 1.780 ;
        RECT  8.760 1.620 10.400 1.780 ;
        RECT  2.230 1.760 3.520 1.920 ;
        RECT  4.160 1.760 5.080 1.920 ;
        RECT  1.340 0.620 1.540 2.100 ;
        RECT  1.140 1.810 1.540 2.100 ;
        RECT  4.920 1.760 5.080 2.100 ;
        RECT  3.360 1.920 4.320 2.080 ;
        RECT  2.230 1.760 2.390 2.100 ;
        RECT  1.140 1.940 2.390 2.100 ;
        RECT  8.080 1.520 8.240 2.100 ;
        RECT  4.920 1.940 8.240 2.100 ;
        RECT  10.560 1.700 11.280 2.100 ;
        RECT  10.960 0.620 11.280 2.100 ;
        RECT  8.760 1.940 11.280 2.100 ;
        RECT  9.600 0.300 11.600 0.460 ;
        RECT  11.440 0.300 11.600 1.230 ;
        RECT  11.440 1.070 12.180 1.230 ;
        RECT  9.600 0.300 9.880 1.460 ;
        LAYER VTPH ;
        RECT  8.750 0.940 10.180 2.400 ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 0.940 ;
        RECT  0.000 0.000 8.750 1.140 ;
        RECT  10.180 0.000 12.800 1.140 ;
    END
END MUX4M1HM

MACRO MUX4M0HM
    CLASS CORE ;
    FOREIGN MUX4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.552  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.010 8.300 1.210 ;
        LAYER ME2 ;
        RECT  8.100 0.840 8.300 1.560 ;
        LAYER ME1 ;
        RECT  8.100 0.860 8.420 1.360 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        ANTENNAGATEAREA 0.154  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.844  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.680 1.010 8.880 1.210 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.880 1.560 ;
        LAYER ME1 ;
        RECT  8.580 0.860 8.920 1.360 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.960 0.440 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.120 3.350 1.280 ;
        RECT  2.500 0.900 2.760 1.280 ;
        RECT  2.440 0.900 2.760 1.100 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.400 1.120 4.900 1.560 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 1.160 7.100 1.440 ;
        RECT  6.100 0.300 6.300 1.440 ;
        RECT  5.120 0.300 6.300 0.460 ;
        RECT  4.360 0.480 5.280 0.640 ;
        RECT  5.120 0.300 5.280 0.640 ;
        RECT  4.360 0.300 4.520 0.640 ;
        RECT  3.600 0.300 4.520 0.460 ;
        RECT  2.920 0.750 3.760 0.950 ;
        RECT  3.600 0.300 3.760 0.950 ;
        RECT  2.920 0.300 3.080 0.950 ;
        RECT  2.460 0.300 3.080 0.730 ;
        RECT  1.020 0.300 3.080 0.460 ;
        RECT  1.020 0.300 1.180 1.580 ;
        END
    END S0
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.220 1.520 12.700 1.820 ;
        RECT  12.500 0.540 12.700 1.820 ;
        RECT  12.220 0.540 12.700 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.640 1.490 11.840 2.540 ;
        RECT  8.400 1.840 8.600 2.540 ;
        RECT  4.480 2.080 4.760 2.540 ;
        RECT  2.920 2.080 3.200 2.540 ;
        RECT  0.140 1.810 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.760 -0.140 11.920 0.880 ;
        RECT  8.400 -0.140 8.600 0.380 ;
        RECT  4.680 -0.140 4.960 0.320 ;
        RECT  3.240 -0.140 3.440 0.560 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.640 0.300 0.840 2.070 ;
        RECT  1.820 0.620 2.300 0.820 ;
        RECT  1.820 0.620 2.020 1.780 ;
        RECT  1.700 1.550 2.020 1.780 ;
        RECT  3.920 0.620 4.200 0.960 ;
        RECT  3.920 0.800 5.280 0.960 ;
        RECT  5.120 0.800 5.280 1.280 ;
        RECT  5.120 1.000 5.600 1.280 ;
        RECT  2.180 1.230 2.340 1.600 ;
        RECT  3.920 0.620 4.080 1.600 ;
        RECT  2.180 1.440 4.080 1.600 ;
        RECT  3.680 1.440 3.960 1.720 ;
        RECT  5.440 0.620 5.920 0.820 ;
        RECT  5.760 0.620 5.920 1.760 ;
        RECT  5.240 1.560 5.920 1.760 ;
        RECT  7.600 0.620 7.920 1.780 ;
        RECT  6.540 0.300 8.240 0.460 ;
        RECT  8.080 0.300 8.240 0.700 ;
        RECT  8.840 0.300 9.280 0.700 ;
        RECT  8.080 0.540 9.280 0.700 ;
        RECT  6.540 0.300 6.820 1.000 ;
        RECT  6.540 0.840 7.420 1.000 ;
        RECT  9.080 0.300 9.280 1.460 ;
        RECT  9.080 1.230 9.360 1.460 ;
        RECT  7.260 0.840 7.420 1.780 ;
        RECT  6.340 1.620 7.420 1.780 ;
        RECT  10.240 0.620 10.800 0.820 ;
        RECT  1.340 0.620 1.620 0.840 ;
        RECT  8.080 1.520 8.920 1.680 ;
        RECT  10.240 0.620 10.400 1.780 ;
        RECT  8.760 1.620 10.400 1.780 ;
        RECT  2.230 1.760 3.520 1.920 ;
        RECT  4.160 1.760 5.080 1.920 ;
        RECT  1.340 0.620 1.540 2.100 ;
        RECT  1.140 1.810 1.540 2.100 ;
        RECT  4.920 1.760 5.080 2.100 ;
        RECT  3.360 1.920 4.320 2.080 ;
        RECT  2.230 1.760 2.390 2.100 ;
        RECT  1.140 1.940 2.390 2.100 ;
        RECT  8.080 1.520 8.240 2.100 ;
        RECT  4.920 1.940 8.240 2.100 ;
        RECT  10.960 0.620 11.280 0.840 ;
        RECT  10.560 1.700 10.840 2.100 ;
        RECT  11.040 0.620 11.280 2.100 ;
        RECT  8.760 1.940 11.280 2.100 ;
        RECT  9.600 0.300 11.600 0.460 ;
        RECT  11.440 0.300 11.600 1.230 ;
        RECT  11.440 1.070 12.180 1.230 ;
        RECT  9.600 0.300 9.880 1.460 ;
        LAYER VTPH ;
        RECT  8.750 0.940 10.180 2.400 ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 0.940 ;
        RECT  0.000 0.000 8.750 1.140 ;
        RECT  10.180 0.000 12.800 1.140 ;
    END
END MUX4M0HM

MACRO MUX3M4HM
    CLASS CORE ;
    FOREIGN MUX3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.454  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.090 1.140 1.290 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.140 1.400 ;
        LAYER ME1 ;
        RECT  0.900 1.020 1.260 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.360 1.120 2.700 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.750 0.840 5.230 1.100 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.560 1.580 1.720 ;
        RECT  1.420 1.300 1.580 1.720 ;
        RECT  0.420 1.130 0.700 1.720 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.188  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.120 3.150 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.900 1.720 6.300 1.920 ;
        RECT  6.100 0.480 6.300 1.920 ;
        RECT  5.900 0.480 6.300 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.460 1.480 6.660 2.540 ;
        RECT  5.440 1.800 5.600 2.540 ;
        RECT  2.540 2.080 2.820 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.460 -0.140 6.660 0.710 ;
        RECT  5.130 -0.140 5.410 0.320 ;
        RECT  2.560 -0.140 2.720 0.640 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.500 0.340 0.860 ;
        RECT  0.100 0.700 2.060 0.860 ;
        RECT  1.900 0.700 2.060 1.420 ;
        RECT  0.100 0.500 0.260 2.080 ;
        RECT  0.100 1.880 0.380 2.080 ;
        RECT  2.880 0.300 3.920 0.460 ;
        RECT  1.540 0.380 2.380 0.540 ;
        RECT  3.720 0.300 3.920 0.640 ;
        RECT  2.220 0.380 2.380 0.960 ;
        RECT  2.880 0.300 3.040 0.960 ;
        RECT  2.220 0.800 3.040 0.960 ;
        RECT  2.000 1.760 3.140 1.920 ;
        RECT  2.980 1.760 3.140 2.100 ;
        RECT  1.500 1.900 2.160 2.060 ;
        RECT  3.790 1.780 3.990 2.100 ;
        RECT  2.980 1.940 3.990 2.100 ;
        RECT  3.200 0.620 3.510 0.820 ;
        RECT  3.310 1.320 4.940 1.520 ;
        RECT  3.310 0.620 3.510 1.780 ;
        RECT  4.240 0.360 4.440 0.640 ;
        RECT  4.240 0.480 5.610 0.640 ;
        RECT  5.450 1.050 5.940 1.250 ;
        RECT  5.450 0.480 5.610 1.640 ;
        RECT  5.120 1.480 5.610 1.640 ;
        RECT  5.120 1.480 5.280 2.020 ;
        RECT  4.340 1.860 5.280 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  2.000 1.140 6.800 2.400 ;
        RECT  0.000 1.220 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
        RECT  0.500 0.000 2.000 1.220 ;
    END
END MUX3M4HM

MACRO MUX3M2HM
    CLASS CORE ;
    FOREIGN MUX3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.090 1.140 1.290 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.140 1.400 ;
        LAYER ME1 ;
        RECT  0.900 1.020 1.260 1.390 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.360 1.120 2.700 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.750 0.840 5.230 1.100 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.550 1.580 1.710 ;
        RECT  1.420 1.300 1.580 1.710 ;
        RECT  0.420 1.130 0.700 1.710 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.120 3.150 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.900 1.720 6.300 1.920 ;
        RECT  6.100 0.480 6.300 1.920 ;
        RECT  5.900 0.480 6.300 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.440 1.800 5.600 2.540 ;
        RECT  2.540 2.080 2.820 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.130 -0.140 5.410 0.320 ;
        RECT  2.560 -0.140 2.720 0.640 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.500 0.340 0.860 ;
        RECT  0.100 0.700 2.060 0.860 ;
        RECT  1.900 0.700 2.060 1.420 ;
        RECT  0.100 0.500 0.260 2.080 ;
        RECT  0.100 1.880 0.380 2.080 ;
        RECT  2.880 0.300 3.920 0.460 ;
        RECT  1.540 0.380 2.380 0.540 ;
        RECT  3.720 0.300 3.920 0.640 ;
        RECT  2.220 0.380 2.380 0.960 ;
        RECT  2.880 0.300 3.040 0.960 ;
        RECT  2.220 0.800 3.040 0.960 ;
        RECT  2.220 1.760 3.140 1.920 ;
        RECT  2.980 1.760 3.140 2.100 ;
        RECT  1.660 1.860 2.380 2.060 ;
        RECT  3.790 1.780 3.990 2.100 ;
        RECT  2.980 1.940 3.990 2.100 ;
        RECT  3.200 0.620 3.510 0.820 ;
        RECT  3.310 1.320 4.940 1.520 ;
        RECT  3.310 0.620 3.510 1.780 ;
        RECT  4.200 0.340 4.480 0.640 ;
        RECT  4.200 0.480 5.610 0.640 ;
        RECT  5.450 1.050 5.840 1.250 ;
        RECT  5.450 0.480 5.610 1.640 ;
        RECT  5.120 1.480 5.610 1.640 ;
        RECT  5.120 1.480 5.280 2.020 ;
        RECT  4.340 1.860 5.280 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  2.000 1.140 6.400 2.400 ;
        RECT  0.000 1.220 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
        RECT  0.500 0.000 2.000 1.220 ;
    END
END MUX3M2HM

MACRO MUX3M1HM
    CLASS CORE ;
    FOREIGN MUX3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.090 1.140 1.290 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.140 1.400 ;
        LAYER ME1 ;
        RECT  0.900 1.020 1.260 1.390 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.360 1.120 2.700 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.750 0.840 5.230 1.100 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.550 1.580 1.710 ;
        RECT  1.420 1.300 1.580 1.710 ;
        RECT  0.420 1.130 0.700 1.710 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.120 3.150 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.900 1.720 6.300 1.920 ;
        RECT  6.100 0.380 6.300 1.920 ;
        RECT  5.900 0.380 6.300 0.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.440 1.800 5.600 2.540 ;
        RECT  2.540 2.080 2.820 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.130 -0.140 5.410 0.320 ;
        RECT  2.560 -0.140 2.720 0.640 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.500 0.340 0.860 ;
        RECT  0.100 0.700 2.060 0.860 ;
        RECT  1.900 0.700 2.060 1.420 ;
        RECT  0.100 0.500 0.260 2.080 ;
        RECT  0.100 1.880 0.380 2.080 ;
        RECT  2.880 0.300 3.920 0.460 ;
        RECT  1.540 0.380 2.380 0.540 ;
        RECT  3.720 0.300 3.920 0.640 ;
        RECT  2.220 0.380 2.380 0.960 ;
        RECT  2.880 0.300 3.040 0.960 ;
        RECT  2.220 0.800 3.040 0.960 ;
        RECT  2.220 1.760 3.140 1.920 ;
        RECT  2.980 1.760 3.140 2.100 ;
        RECT  1.660 1.860 2.380 2.060 ;
        RECT  3.790 1.780 3.990 2.100 ;
        RECT  2.980 1.940 3.990 2.100 ;
        RECT  3.200 0.620 3.510 0.820 ;
        RECT  3.310 1.320 4.940 1.520 ;
        RECT  3.310 0.620 3.510 1.780 ;
        RECT  4.200 0.340 4.480 0.640 ;
        RECT  4.200 0.480 5.610 0.640 ;
        RECT  5.450 1.050 5.840 1.250 ;
        RECT  5.450 0.480 5.610 1.640 ;
        RECT  5.120 1.480 5.610 1.640 ;
        RECT  5.120 1.480 5.280 2.020 ;
        RECT  4.340 1.860 5.280 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  2.000 1.140 6.400 2.400 ;
        RECT  0.000 1.220 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
        RECT  0.500 0.000 2.000 1.220 ;
    END
END MUX3M1HM

MACRO MUX3M0HM
    CLASS CORE ;
    FOREIGN MUX3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.090 1.140 1.290 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.140 1.400 ;
        LAYER ME1 ;
        RECT  0.900 1.020 1.260 1.390 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.360 1.120 2.700 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.750 0.840 5.230 1.100 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.550 1.580 1.710 ;
        RECT  1.420 1.300 1.580 1.710 ;
        RECT  0.420 1.130 0.700 1.710 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.120 3.150 1.560 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.900 1.800 6.300 2.000 ;
        RECT  6.100 0.340 6.300 2.000 ;
        RECT  5.900 0.340 6.300 0.540 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.440 1.800 5.600 2.540 ;
        RECT  2.540 2.080 2.820 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.130 -0.140 5.410 0.320 ;
        RECT  2.560 -0.140 2.720 0.640 ;
        RECT  0.660 -0.140 0.940 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.500 0.340 0.860 ;
        RECT  0.100 0.700 2.060 0.860 ;
        RECT  1.900 0.700 2.060 1.420 ;
        RECT  0.100 0.500 0.260 2.080 ;
        RECT  0.100 1.880 0.380 2.080 ;
        RECT  2.880 0.300 3.920 0.460 ;
        RECT  1.540 0.380 2.380 0.540 ;
        RECT  3.720 0.300 3.920 0.640 ;
        RECT  2.220 0.380 2.380 0.960 ;
        RECT  2.880 0.300 3.040 0.960 ;
        RECT  2.220 0.800 3.040 0.960 ;
        RECT  2.220 1.760 3.140 1.920 ;
        RECT  2.980 1.760 3.140 2.100 ;
        RECT  1.660 1.860 2.380 2.060 ;
        RECT  3.790 1.780 3.990 2.100 ;
        RECT  2.980 1.940 3.990 2.100 ;
        RECT  3.200 0.620 3.510 0.820 ;
        RECT  3.310 1.320 4.940 1.520 ;
        RECT  3.310 0.620 3.510 1.780 ;
        RECT  4.200 0.340 4.480 0.640 ;
        RECT  4.200 0.480 5.680 0.640 ;
        RECT  5.520 0.480 5.680 1.640 ;
        RECT  5.120 1.480 5.680 1.640 ;
        RECT  5.120 1.480 5.280 2.020 ;
        RECT  4.340 1.860 5.280 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  2.000 1.140 6.400 2.400 ;
        RECT  0.000 1.220 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
        RECT  0.500 0.000 2.000 1.220 ;
    END
END MUX3M0HM

MACRO MUX2M8HM
    CLASS CORE ;
    FOREIGN MUX2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.620 1.060 3.900 1.660 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.820 1.300 1.340 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.209  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.300 2.090 1.180 ;
        RECT  1.100 0.300 2.090 0.460 ;
        RECT  0.500 0.500 1.300 0.660 ;
        RECT  1.100 0.300 1.300 0.660 ;
        RECT  0.500 0.500 0.740 1.340 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.500 0.390 5.780 2.080 ;
        RECT  4.480 0.880 5.780 1.160 ;
        RECT  4.480 0.390 4.740 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  6.020 1.440 6.300 2.540 ;
        RECT  4.980 1.440 5.260 2.540 ;
        RECT  3.960 1.820 4.220 2.540 ;
        RECT  0.660 1.880 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  6.020 -0.140 6.300 0.560 ;
        RECT  4.980 -0.140 5.260 0.560 ;
        RECT  3.960 -0.140 4.220 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.620 1.740 1.720 ;
        RECT  2.820 1.010 3.100 1.290 ;
        RECT  0.100 0.310 0.340 1.720 ;
        RECT  0.100 1.500 1.300 1.720 ;
        RECT  1.110 1.500 1.300 2.100 ;
        RECT  2.820 1.010 3.040 2.100 ;
        RECT  1.110 1.940 3.040 2.100 ;
        RECT  3.160 0.620 3.460 0.840 ;
        RECT  3.260 0.620 3.460 2.080 ;
        RECT  3.200 1.440 3.460 2.080 ;
        RECT  2.250 0.300 3.800 0.460 ;
        RECT  3.640 0.300 3.800 0.880 ;
        RECT  3.640 0.720 4.320 0.880 ;
        RECT  4.060 0.720 4.320 1.290 ;
        RECT  2.250 0.300 2.500 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END MUX2M8HM

MACRO MUX2M6HM
    CLASS CORE ;
    FOREIGN MUX2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.060 2.880 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.180  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.060 1.940 2.260 2.100 ;
        RECT  2.100 0.700 2.260 2.100 ;
        RECT  1.060 1.480 1.220 2.100 ;
        RECT  0.500 1.480 1.220 1.640 ;
        RECT  0.500 1.010 0.700 1.640 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.420 0.430 4.620 2.100 ;
        RECT  3.540 0.900 4.620 1.100 ;
        RECT  3.340 1.520 3.700 2.080 ;
        RECT  3.540 0.320 3.700 2.080 ;
        RECT  3.340 0.320 3.700 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.900 1.480 4.100 2.540 ;
        RECT  2.860 1.840 3.060 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.900 -0.140 4.100 0.710 ;
        RECT  2.860 -0.140 3.060 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.520 1.620 0.680 ;
        RECT  1.420 0.520 1.620 1.180 ;
        RECT  0.140 0.520 0.340 1.740 ;
        RECT  1.780 0.320 2.660 0.520 ;
        RECT  2.500 0.320 2.660 0.880 ;
        RECT  2.500 0.720 3.380 0.880 ;
        RECT  3.220 0.720 3.380 1.330 ;
        RECT  1.780 0.320 1.940 1.680 ;
        RECT  1.540 1.480 1.940 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END MUX2M6HM

MACRO MUX2M4HM
    CLASS CORE ;
    FOREIGN MUX2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.060 2.880 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.180  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.060 1.940 2.260 2.100 ;
        RECT  2.100 0.700 2.260 2.100 ;
        RECT  1.060 1.480 1.220 2.100 ;
        RECT  0.500 1.480 1.220 1.640 ;
        RECT  0.500 1.010 0.700 1.640 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.520 3.700 2.080 ;
        RECT  3.540 0.320 3.700 2.080 ;
        RECT  3.340 0.320 3.700 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.900 1.480 4.100 2.540 ;
        RECT  2.860 1.840 3.060 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.900 -0.140 4.100 0.710 ;
        RECT  2.860 -0.140 3.060 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.500 1.480 0.660 ;
        RECT  1.320 0.500 1.480 1.180 ;
        RECT  1.320 0.900 1.620 1.180 ;
        RECT  0.140 0.500 0.340 1.740 ;
        RECT  1.780 0.320 2.660 0.520 ;
        RECT  2.500 0.320 2.660 0.880 ;
        RECT  2.500 0.720 3.380 0.880 ;
        RECT  3.220 0.720 3.380 1.330 ;
        RECT  1.780 0.320 1.940 1.680 ;
        RECT  1.540 1.480 1.940 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MUX2M4HM

MACRO MUX2M3HM
    CLASS CORE ;
    FOREIGN MUX2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.097  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.090 2.910 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.166  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.060 1.940 2.260 2.100 ;
        RECT  2.100 0.700 2.260 2.100 ;
        RECT  1.060 1.480 1.220 2.100 ;
        RECT  0.500 1.480 1.220 1.640 ;
        RECT  0.500 1.010 0.700 1.640 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.372  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.390 1.620 3.900 1.820 ;
        RECT  3.700 0.320 3.900 1.820 ;
        RECT  3.390 0.320 3.900 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.060 1.580 4.260 2.540 ;
        RECT  2.870 1.760 3.150 2.540 ;
        RECT  0.700 1.800 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.620 ;
        RECT  2.910 -0.140 3.110 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.480 1.480 0.640 ;
        RECT  1.320 0.480 1.480 1.180 ;
        RECT  1.320 0.900 1.620 1.180 ;
        RECT  0.140 0.390 0.340 1.980 ;
        RECT  1.780 0.320 2.710 0.520 ;
        RECT  2.550 0.320 2.710 0.880 ;
        RECT  2.550 0.720 3.430 0.880 ;
        RECT  3.270 0.720 3.430 1.330 ;
        RECT  1.780 0.320 1.940 1.680 ;
        RECT  1.540 1.480 1.940 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MUX2M3HM

MACRO MUX2M2HM
    CLASS CORE ;
    FOREIGN MUX2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.060 2.700 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 0.700 2.160 0.900 ;
        RECT  0.500 1.520 1.940 1.680 ;
        RECT  1.780 0.700 1.940 1.680 ;
        RECT  0.500 1.010 0.700 1.680 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.521  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.390 3.500 2.080 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.640 -0.140 2.840 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.580 2.080 2.860 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.480 0.680 ;
        RECT  1.320 0.480 1.480 1.260 ;
        RECT  1.320 0.980 1.620 1.260 ;
        RECT  0.100 0.480 0.300 2.080 ;
        RECT  0.100 1.880 0.390 2.080 ;
        RECT  1.660 0.340 2.480 0.500 ;
        RECT  2.320 0.340 2.480 0.880 ;
        RECT  2.320 0.720 3.060 0.880 ;
        RECT  2.900 0.720 3.060 1.880 ;
        RECT  2.100 1.720 3.060 1.880 ;
        RECT  2.100 1.720 2.260 2.060 ;
        RECT  1.420 1.900 2.260 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MUX2M2HM

MACRO MUX2M1HM
    CLASS CORE ;
    FOREIGN MUX2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.160 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.060 2.700 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 0.700 2.160 0.900 ;
        RECT  0.500 1.520 1.940 1.680 ;
        RECT  1.780 0.700 1.940 1.680 ;
        RECT  0.500 1.010 0.700 1.680 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.365  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.390 3.500 1.850 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.640 -0.140 2.840 0.560 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.580 2.080 2.860 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.480 0.680 ;
        RECT  1.320 0.480 1.480 1.260 ;
        RECT  1.320 0.980 1.620 1.260 ;
        RECT  0.100 0.480 0.300 2.080 ;
        RECT  0.100 1.880 0.390 2.080 ;
        RECT  1.660 0.340 2.480 0.500 ;
        RECT  2.320 0.340 2.480 0.880 ;
        RECT  2.320 0.720 3.060 0.880 ;
        RECT  2.900 0.720 3.060 1.880 ;
        RECT  2.100 1.720 3.060 1.880 ;
        RECT  2.100 1.720 2.260 2.060 ;
        RECT  1.420 1.900 2.260 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MUX2M1HM

MACRO MUX2M0HM
    CLASS CORE ;
    FOREIGN MUX2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.620 1.060 3.900 1.660 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.820 1.300 1.340 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.113  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.940 0.300 2.130 1.180 ;
        RECT  1.140 0.300 2.130 0.460 ;
        RECT  0.500 0.500 1.300 0.660 ;
        RECT  1.140 0.300 1.300 0.660 ;
        RECT  0.500 0.500 0.740 1.340 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.440 0.300 4.700 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.920 1.820 4.180 2.540 ;
        RECT  0.700 1.880 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.500 0.620 1.780 1.720 ;
        RECT  2.820 1.010 3.100 1.290 ;
        RECT  0.100 0.310 0.340 1.720 ;
        RECT  0.100 1.500 1.340 1.720 ;
        RECT  1.150 1.500 1.340 2.100 ;
        RECT  2.820 1.010 3.040 2.100 ;
        RECT  1.150 1.940 3.040 2.100 ;
        RECT  3.160 0.620 3.460 0.840 ;
        RECT  3.260 0.620 3.460 1.780 ;
        RECT  3.200 1.500 3.460 1.780 ;
        RECT  2.330 0.300 3.780 0.460 ;
        RECT  3.620 0.300 3.780 0.880 ;
        RECT  3.620 0.720 4.280 0.880 ;
        RECT  4.060 0.720 4.280 1.290 ;
        RECT  2.330 0.300 2.550 1.780 ;
        RECT  2.190 1.500 2.550 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END MUX2M0HM

MACRO MOAI22M4HM
    CLASS CORE ;
    FOREIGN MOAI22M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.420 1.290 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 0.900 1.160 1.290 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 2.040 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 0.840 2.700 1.260 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.500 1.460 4.300 1.740 ;
        RECT  4.100 0.680 4.300 1.740 ;
        RECT  3.500 0.680 4.300 0.860 ;
        RECT  3.500 0.390 3.780 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.900 4.300 2.540 ;
        RECT  2.980 1.840 3.260 2.540 ;
        RECT  0.100 2.020 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.020 -0.140 4.300 0.520 ;
        RECT  2.540 -0.140 3.220 0.320 ;
        RECT  1.100 -0.140 1.380 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.520 1.500 0.740 ;
        RECT  1.340 0.520 1.500 1.700 ;
        RECT  0.100 1.490 1.500 1.700 ;
        RECT  1.460 1.860 2.780 2.080 ;
        RECT  1.660 0.410 1.940 0.680 ;
        RECT  1.660 0.520 3.300 0.680 ;
        RECT  3.100 1.020 3.900 1.300 ;
        RECT  3.100 0.520 3.300 1.660 ;
        RECT  1.980 1.440 3.300 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MOAI22M4HM

MACRO MOAI22M2HM
    CLASS CORE ;
    FOREIGN MOAI22M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.080 2.200 1.340 ;
        RECT  1.700 0.840 1.960 1.340 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.040 2.700 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.420 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.220 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.650 1.730 3.100 1.890 ;
        RECT  2.900 0.720 3.100 1.890 ;
        RECT  2.220 0.720 3.100 0.880 ;
        RECT  2.220 0.620 2.540 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.580 2.050 2.860 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        RECT  0.100 2.080 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.100 -0.140 1.380 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.560 0.420 0.880 ;
        RECT  0.140 0.720 1.540 0.880 ;
        RECT  1.380 0.720 1.540 1.290 ;
        RECT  0.580 0.720 0.740 1.950 ;
        RECT  0.580 1.730 0.900 1.950 ;
        RECT  1.700 0.300 3.020 0.460 ;
        RECT  2.740 0.300 3.020 0.560 ;
        RECT  1.700 0.300 1.980 0.620 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MOAI22M2HM

MACRO MOAI22M1HM
    CLASS CORE ;
    FOREIGN MOAI22M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 2.100 1.340 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.400 1.040 2.700 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.420 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.220 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.366  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.730 3.100 1.890 ;
        RECT  2.900 0.720 3.100 1.890 ;
        RECT  2.260 0.720 3.100 0.880 ;
        RECT  2.260 0.620 2.540 0.880 ;
        RECT  1.700 1.600 1.980 1.890 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.580 2.050 2.860 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        RECT  0.100 2.080 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.100 -0.140 1.380 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.410 0.420 0.880 ;
        RECT  0.140 0.720 1.540 0.880 ;
        RECT  1.380 0.720 1.540 1.290 ;
        RECT  0.580 0.720 0.740 2.010 ;
        RECT  0.580 1.730 0.900 2.010 ;
        RECT  1.720 0.300 3.100 0.460 ;
        RECT  2.820 0.300 3.100 0.560 ;
        RECT  1.720 0.300 1.940 0.620 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MOAI22M1HM

MACRO MOAI22M0HM
    CLASS CORE ;
    FOREIGN MOAI22M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 2.100 1.340 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.110 2.720 1.560 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.420 1.560 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.160 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.345  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.740 1.730 3.100 1.890 ;
        RECT  2.900 0.790 3.100 1.890 ;
        RECT  2.260 0.790 3.100 0.950 ;
        RECT  2.260 0.620 2.540 0.950 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.660 2.050 2.940 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        RECT  0.100 2.080 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.060 -0.140 1.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.410 0.420 0.880 ;
        RECT  0.140 0.720 1.540 0.880 ;
        RECT  1.320 0.720 1.540 1.250 ;
        RECT  0.580 0.720 0.740 2.010 ;
        RECT  0.580 1.730 0.900 2.010 ;
        RECT  1.660 0.300 3.100 0.460 ;
        RECT  1.660 0.300 1.940 0.520 ;
        RECT  2.820 0.300 3.100 0.630 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MOAI22M0HM

MACRO MAOI22M4HM
    CLASS CORE ;
    FOREIGN MAOI22M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.011  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.700 1.080 2.200 1.400 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.864  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.140 2.700 1.340 ;
        LAYER ME2 ;
        RECT  2.500 1.040 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.040 2.860 1.420 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 0.600 1.400 ;
        RECT  0.100 1.080 0.300 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.040 1.180 1.540 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.460 1.580 4.300 1.740 ;
        RECT  4.100 0.680 4.300 1.740 ;
        RECT  3.540 0.680 4.300 0.880 ;
        RECT  3.540 0.410 3.740 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.900 4.300 2.540 ;
        RECT  2.980 1.900 3.260 2.540 ;
        RECT  2.500 1.900 2.780 2.540 ;
        RECT  1.100 2.080 1.380 2.540 ;
        RECT  0.100 2.080 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.020 -0.140 4.300 0.520 ;
        RECT  2.980 -0.140 3.260 0.520 ;
        RECT  0.940 -0.140 1.140 0.400 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.520 0.320 0.880 ;
        RECT  0.160 0.720 1.500 0.880 ;
        RECT  1.340 0.720 1.500 1.860 ;
        RECT  0.540 1.700 1.500 1.860 ;
        RECT  1.460 0.300 2.780 0.460 ;
        RECT  1.460 0.300 1.740 0.560 ;
        RECT  2.500 0.300 2.780 0.560 ;
        RECT  1.980 0.620 2.260 0.880 ;
        RECT  1.980 0.720 3.300 0.880 ;
        RECT  3.100 1.060 3.900 1.340 ;
        RECT  3.100 0.720 3.300 1.740 ;
        RECT  1.700 1.580 3.300 1.740 ;
        RECT  1.700 1.580 1.900 2.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MAOI22M4HM

MACRO MAOI22M2HM
    CLASS CORE ;
    FOREIGN MAOI22M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.020 2.160 1.300 ;
        RECT  1.700 1.020 1.900 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.840 2.740 1.370 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.420 1.330 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.120 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.452  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.180 1.560 3.100 1.720 ;
        RECT  2.900 0.520 3.100 1.720 ;
        RECT  1.660 0.520 3.100 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.100 2.080 1.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  1.180 -0.140 1.380 0.400 ;
        RECT  0.140 -0.140 0.340 0.400 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.620 0.940 0.780 ;
        RECT  0.580 0.620 0.740 1.920 ;
        RECT  1.380 1.010 1.540 1.920 ;
        RECT  0.180 1.760 1.540 1.920 ;
        RECT  0.180 1.760 0.460 2.060 ;
        RECT  1.700 1.900 3.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MAOI22M2HM

MACRO MAOI22M1HM
    CLASS CORE ;
    FOREIGN MAOI22M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.020 2.160 1.300 ;
        RECT  1.700 1.020 1.900 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.840 2.740 1.400 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.420 1.330 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.120 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.469  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.110 1.580 3.100 1.740 ;
        RECT  2.900 0.520 3.100 1.740 ;
        RECT  1.700 0.520 3.100 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  0.980 1.880 1.260 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        RECT  1.180 -0.140 1.380 0.400 ;
        RECT  0.140 -0.140 0.340 0.400 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.620 1.540 0.780 ;
        RECT  1.380 0.620 1.540 1.370 ;
        RECT  0.580 0.620 0.740 2.060 ;
        RECT  0.100 1.860 0.740 2.060 ;
        RECT  1.540 1.900 3.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MAOI22M1HM

MACRO MAOI22M0HM
    CLASS CORE ;
    FOREIGN MAOI22M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.020 2.160 1.300 ;
        RECT  1.700 1.020 1.900 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.840 2.740 1.400 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.420 1.330 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.120 1.560 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.429  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.110 1.580 3.100 1.740 ;
        RECT  2.900 0.520 3.100 1.740 ;
        RECT  1.700 0.520 3.100 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  0.980 1.900 1.260 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        RECT  1.180 -0.140 1.380 0.400 ;
        RECT  0.140 -0.140 0.340 0.400 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 0.620 1.540 0.780 ;
        RECT  1.380 0.620 1.540 1.370 ;
        RECT  0.580 0.620 0.740 2.060 ;
        RECT  0.100 1.840 0.740 2.060 ;
        RECT  1.540 1.900 3.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MAOI22M0HM

MACRO MAOI222M4HM
    CLASS CORE ;
    FOREIGN MAOI222M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.058  LAYER ME1  ;
        ANTENNAGATEAREA 0.058  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.222  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.150 1.900 1.350 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.500 1.060 1.940 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.540 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.580 2.340 1.740 ;
        RECT  2.100 1.080 2.340 1.740 ;
        RECT  1.140 1.100 1.340 1.740 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.400 1.510 5.100 1.710 ;
        RECT  4.900 0.680 5.100 1.710 ;
        RECT  4.400 0.680 5.100 0.880 ;
        RECT  4.400 1.510 4.600 2.100 ;
        RECT  4.400 0.410 4.600 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  4.860 1.900 5.140 2.540 ;
        RECT  3.820 1.900 4.100 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  4.860 -0.140 5.140 0.520 ;
        RECT  3.820 -0.140 4.100 0.520 ;
        RECT  1.900 -0.140 2.180 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 1.580 0.460 ;
        RECT  1.300 0.300 1.580 0.540 ;
        RECT  0.100 0.300 0.380 0.780 ;
        RECT  0.100 1.900 1.620 2.100 ;
        RECT  0.700 0.700 3.100 0.900 ;
        RECT  2.820 1.080 3.760 1.280 ;
        RECT  0.700 0.620 0.980 1.740 ;
        RECT  2.820 0.560 3.100 2.080 ;
        RECT  3.350 0.300 3.530 0.870 ;
        RECT  3.350 0.690 4.240 0.870 ;
        RECT  4.060 1.040 4.740 1.320 ;
        RECT  4.060 0.690 4.240 1.600 ;
        RECT  3.360 1.440 4.240 1.600 ;
        RECT  3.360 1.440 3.560 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END MAOI222M4HM

MACRO MAOI222M2HM
    CLASS CORE ;
    FOREIGN MAOI222M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.640 0.980 1.920 1.140 ;
        RECT  0.640 0.440 0.800 1.140 ;
        RECT  0.500 0.440 0.800 0.760 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.180 1.300 2.340 1.460 ;
        RECT  2.180 1.020 2.340 1.460 ;
        RECT  0.500 1.300 0.700 1.960 ;
        RECT  0.180 1.300 0.700 1.480 ;
        RECT  0.180 1.120 0.460 1.480 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.060 0.840 3.500 1.310 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.620 2.700 1.780 ;
        RECT  2.500 0.620 2.700 1.780 ;
        RECT  0.960 0.620 2.700 0.780 ;
        RECT  0.960 0.380 1.200 0.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.180 1.480 3.400 2.540 ;
        RECT  0.140 1.690 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.250 -0.140 3.410 0.650 ;
        RECT  0.160 -0.140 0.320 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.380 1.940 2.940 2.100 ;
        RECT  1.380 0.300 2.940 0.460 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MAOI222M2HM

MACRO MAOI222M1HM
    CLASS CORE ;
    FOREIGN MAOI222M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.640 0.980 1.920 1.140 ;
        RECT  0.640 0.440 0.800 1.140 ;
        RECT  0.500 0.440 0.800 0.760 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.180 1.300 2.340 1.460 ;
        RECT  2.120 1.020 2.340 1.460 ;
        RECT  0.500 1.300 0.700 1.960 ;
        RECT  0.180 1.300 0.700 1.480 ;
        RECT  0.180 1.210 0.460 1.480 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.060 0.840 3.500 1.310 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.739  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.620 2.700 1.780 ;
        RECT  2.500 0.620 2.700 1.780 ;
        RECT  0.960 0.620 2.700 0.780 ;
        RECT  0.960 0.320 1.200 0.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.240 1.580 3.400 2.540 ;
        RECT  0.140 1.690 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.250 -0.140 3.410 0.650 ;
        RECT  0.160 -0.140 0.320 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.380 1.940 2.940 2.100 ;
        RECT  1.380 0.300 2.940 0.460 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MAOI222M1HM

MACRO MAOI222M0HM
    CLASS CORE ;
    FOREIGN MAOI222M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.520 1.350 2.800 1.630 ;
        RECT  1.710 1.700 2.680 1.920 ;
        RECT  2.520 1.350 2.680 1.920 ;
        RECT  1.220 1.580 1.870 1.740 ;
        RECT  1.220 1.260 1.380 1.740 ;
        RECT  0.540 1.260 1.380 1.420 ;
        RECT  0.540 1.000 0.760 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.160 0.940 2.760 1.100 ;
        RECT  2.120 0.800 2.760 1.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.260 2.360 1.500 ;
        RECT  1.640 1.260 2.360 1.420 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.721  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 1.820 3.120 2.100 ;
        RECT  2.960 0.300 3.120 2.100 ;
        RECT  2.820 0.300 3.120 0.640 ;
        RECT  1.780 0.480 3.120 0.640 ;
        RECT  0.700 0.620 1.940 0.780 ;
        RECT  0.100 1.580 1.020 1.740 ;
        RECT  0.100 0.680 0.980 0.840 ;
        RECT  0.100 0.680 0.300 1.740 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  1.900 -0.140 2.180 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.900 1.540 2.100 ;
        RECT  0.100 0.300 1.620 0.460 ;
        RECT  0.100 0.300 0.380 0.520 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END MAOI222M0HM

MACRO MAOI2223M4HM
    CLASS CORE ;
    FOREIGN MAOI2223M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.190 2.620 1.620 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.800 2.320 0.960 ;
        RECT  0.100 0.800 0.300 1.160 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 1.790 1.280 ;
        RECT  0.500 1.120 0.700 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.048  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.840 3.500 1.370 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.500 1.510 6.300 1.710 ;
        RECT  6.100 0.700 6.300 1.710 ;
        RECT  5.510 0.700 6.300 0.900 ;
        RECT  5.500 1.510 5.780 2.100 ;
        RECT  5.510 0.380 5.760 0.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  6.020 1.900 6.300 2.540 ;
        RECT  4.980 1.900 5.260 2.540 ;
        RECT  3.980 1.900 4.260 2.540 ;
        RECT  1.300 1.900 1.580 2.540 ;
        RECT  0.100 1.920 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  6.020 -0.140 6.300 0.540 ;
        RECT  4.980 -0.140 5.260 0.540 ;
        RECT  3.980 -0.140 4.260 0.760 ;
        RECT  1.300 -0.140 1.580 0.320 ;
        RECT  0.100 -0.140 0.380 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.760 0.300 3.660 0.460 ;
        RECT  1.760 0.300 1.920 0.640 ;
        RECT  0.660 0.480 1.920 0.640 ;
        RECT  3.380 0.300 3.660 0.680 ;
        RECT  0.960 1.580 1.900 1.740 ;
        RECT  1.740 1.580 1.900 2.060 ;
        RECT  0.660 1.740 1.120 1.900 ;
        RECT  1.740 1.900 3.700 2.060 ;
        RECT  2.700 0.620 3.060 0.880 ;
        RECT  4.100 1.200 4.920 1.420 ;
        RECT  2.780 0.620 3.060 1.740 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  2.780 1.580 4.300 1.740 ;
        RECT  4.460 0.340 4.740 1.010 ;
        RECT  4.460 0.830 5.260 1.010 ;
        RECT  5.080 1.060 5.900 1.340 ;
        RECT  5.080 0.830 5.260 1.740 ;
        RECT  4.510 1.580 5.260 1.740 ;
        RECT  4.510 1.580 4.690 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END MAOI2223M4HM

MACRO MAOI2223M2HM
    CLASS CORE ;
    FOREIGN MAOI2223M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.900 3.780 1.140 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.265  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.300 4.300 1.460 ;
        RECT  4.080 0.840 4.300 1.460 ;
        RECT  2.860 1.020 3.020 1.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.265  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.440 2.340 1.600 ;
        RECT  2.180 1.020 2.340 1.600 ;
        RECT  0.100 1.080 0.340 1.600 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.265  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 1.960 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.640  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.620 3.180 1.780 ;
        RECT  2.500 0.620 3.100 0.820 ;
        RECT  2.500 0.620 2.700 1.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.000 1.840 4.240 2.540 ;
        RECT  1.420 2.080 1.700 2.540 ;
        RECT  0.380 1.840 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.980 -0.140 4.260 0.500 ;
        RECT  1.480 -0.140 1.640 0.600 ;
        RECT  0.380 -0.140 0.580 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 1.760 2.060 1.920 ;
        RECT  1.900 1.760 2.060 2.100 ;
        RECT  3.460 1.900 3.740 2.100 ;
        RECT  1.900 1.940 3.740 2.100 ;
        RECT  1.800 0.300 3.770 0.460 ;
        RECT  3.460 0.300 3.770 0.500 ;
        RECT  0.920 0.300 1.080 0.920 ;
        RECT  1.800 0.300 1.960 0.920 ;
        RECT  0.920 0.760 1.960 0.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MAOI2223M2HM

MACRO MAOI2223M1HM
    CLASS CORE ;
    FOREIGN MAOI2223M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.088  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.900 3.700 1.140 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.187  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.300 4.300 1.460 ;
        RECT  4.080 0.840 4.300 1.460 ;
        RECT  2.860 1.020 3.020 1.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.187  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.440 2.340 1.600 ;
        RECT  2.180 1.020 2.340 1.600 ;
        RECT  0.100 1.080 0.340 1.600 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.187  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 1.960 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.509  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.620 3.180 1.780 ;
        RECT  2.500 0.620 3.100 0.820 ;
        RECT  2.500 0.620 2.700 1.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.000 1.760 4.240 2.540 ;
        RECT  1.420 2.080 1.700 2.540 ;
        RECT  0.380 1.760 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.980 -0.140 4.260 0.500 ;
        RECT  1.480 -0.140 1.640 0.600 ;
        RECT  0.380 -0.140 0.580 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.820 1.760 2.060 1.920 ;
        RECT  1.900 1.760 2.060 2.100 ;
        RECT  3.460 1.820 3.740 2.100 ;
        RECT  1.900 1.940 3.740 2.100 ;
        RECT  1.800 0.300 3.770 0.460 ;
        RECT  3.460 0.300 3.770 0.500 ;
        RECT  0.880 0.300 1.120 0.920 ;
        RECT  1.800 0.300 1.960 0.920 ;
        RECT  0.880 0.760 1.960 0.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MAOI2223M1HM

MACRO MAOI2223M0HM
    CLASS CORE ;
    FOREIGN MAOI2223M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.780 1.300 4.300 1.460 ;
        RECT  4.080 0.840 4.300 1.460 ;
        RECT  2.780 1.100 2.940 1.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.440 2.280 1.600 ;
        RECT  2.000 1.340 2.280 1.600 ;
        RECT  0.100 1.080 0.340 1.600 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 1.840 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.240 0.660 3.580 1.140 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.512  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.620 3.180 1.780 ;
        RECT  2.440 0.620 3.050 0.780 ;
        RECT  2.440 0.620 2.600 1.780 ;
        RECT  2.040 0.900 2.600 1.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.000 1.760 4.240 2.540 ;
        RECT  1.300 2.080 1.580 2.540 ;
        RECT  0.100 1.760 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.020 -0.140 4.300 0.500 ;
        RECT  1.380 -0.140 1.540 0.600 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.720 0.300 3.700 0.460 ;
        RECT  0.660 0.340 1.220 0.500 ;
        RECT  3.420 0.300 3.700 0.500 ;
        RECT  1.060 0.340 1.220 0.920 ;
        RECT  1.720 0.300 1.880 0.920 ;
        RECT  1.060 0.760 1.880 0.920 ;
        RECT  0.680 1.760 2.060 1.920 ;
        RECT  1.900 1.760 2.060 2.100 ;
        RECT  3.460 1.820 3.740 2.100 ;
        RECT  1.900 1.940 3.740 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MAOI2223M0HM

MACRO MAO222M4HM
    CLASS CORE ;
    FOREIGN MAO222M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.280  LAYER ME1  ;
        ANTENNAGATEAREA 0.280  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.691  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.160 2.300 1.360 ;
        LAYER ME2 ;
        RECT  2.100 0.900 2.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.260 2.560 1.420 ;
        RECT  2.000 1.120 2.560 1.420 ;
        RECT  0.100 0.960 0.320 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.650  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.830 1.170 3.030 1.370 ;
        LAYER ME2 ;
        RECT  2.830 0.900 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.720 1.120 3.160 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.280  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.820 0.980 1.100 ;
        RECT  0.500 0.440 0.700 1.100 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.650 1.510 4.300 1.740 ;
        RECT  4.100 0.660 4.300 1.740 ;
        RECT  3.650 0.660 4.300 0.820 ;
        RECT  3.500 1.900 3.850 2.100 ;
        RECT  3.650 1.510 3.850 2.100 ;
        RECT  3.650 0.300 3.850 0.820 ;
        RECT  3.500 0.300 3.850 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.900 4.300 2.540 ;
        RECT  2.980 1.900 3.260 2.540 ;
        RECT  0.100 1.840 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.020 -0.140 4.300 0.500 ;
        RECT  2.980 -0.140 3.260 0.500 ;
        RECT  0.100 -0.140 0.320 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.480 0.300 2.740 0.460 ;
        RECT  2.460 0.300 2.740 0.540 ;
        RECT  1.480 0.300 1.700 0.600 ;
        RECT  1.380 1.900 2.780 2.100 ;
        RECT  0.890 0.300 1.320 0.620 ;
        RECT  1.160 0.300 1.320 0.960 ;
        RECT  1.940 0.620 2.220 0.960 ;
        RECT  1.160 0.760 3.490 0.960 ;
        RECT  3.320 1.020 3.940 1.300 ;
        RECT  3.320 0.760 3.490 1.740 ;
        RECT  0.940 1.580 3.490 1.740 ;
        RECT  0.940 1.580 1.220 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END MAO222M4HM

MACRO MAO222M2HM
    CLASS CORE ;
    FOREIGN MAO222M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.160 1.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 1.260 2.700 1.420 ;
        RECT  2.460 0.840 2.700 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.900 1.960 1.100 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.420 3.500 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.620 -0.140 2.900 0.340 ;
        RECT  0.580 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 1.580 1.540 1.740 ;
        RECT  0.160 1.580 0.320 1.940 ;
        RECT  1.720 0.300 1.880 0.660 ;
        RECT  1.720 0.500 3.100 0.660 ;
        RECT  2.940 0.500 3.100 1.740 ;
        RECT  1.700 1.580 3.100 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MAO222M2HM

MACRO MAO222M1HM
    CLASS CORE ;
    FOREIGN MAO222M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.160 1.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 1.260 2.700 1.420 ;
        RECT  2.460 0.840 2.700 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.900 1.960 1.100 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.313  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.450 3.500 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.620 -0.140 2.900 0.340 ;
        RECT  0.580 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 1.580 1.540 1.740 ;
        RECT  0.160 1.580 0.320 1.940 ;
        RECT  1.720 0.300 1.880 0.660 ;
        RECT  1.720 0.500 3.100 0.660 ;
        RECT  2.940 0.500 3.100 1.740 ;
        RECT  1.700 1.580 3.100 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MAO222M1HM

MACRO MAO222M0HM
    CLASS CORE ;
    FOREIGN MAO222M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.160 1.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 1.260 2.700 1.420 ;
        RECT  2.460 0.840 2.700 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.440 0.900 1.960 1.100 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.241  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.500 3.500 1.770 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.620 -0.140 2.900 0.340 ;
        RECT  0.580 -0.140 0.860 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 1.580 1.540 1.740 ;
        RECT  0.160 1.580 0.320 1.940 ;
        RECT  1.720 0.300 1.880 0.660 ;
        RECT  1.720 0.500 3.100 0.660 ;
        RECT  2.940 0.500 3.100 1.740 ;
        RECT  1.700 1.580 3.100 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END MAO222M0HM

MACRO LARSM4HM
    CLASS CORE ;
    FOREIGN LARSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.454  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.500 0.760 1.700 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.660 1.700 1.160 ;
        LAYER ME1 ;
        RECT  1.400 0.700 1.880 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.140 1.280 ;
        RECT  2.060 1.080 3.140 1.280 ;
        RECT  2.060 0.960 2.340 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.640 0.390 7.900 2.080 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.480 0.430 6.760 1.600 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.080 3.960 1.280 ;
        RECT  3.300 0.640 3.500 1.280 ;
        RECT  2.040 0.640 3.500 0.800 ;
        RECT  2.040 0.320 2.200 0.800 ;
        RECT  1.040 0.320 2.200 0.480 ;
        RECT  1.040 0.320 1.240 0.940 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.760 5.180 1.160 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.160 1.480 8.360 2.540 ;
        RECT  7.040 2.080 7.320 2.540 ;
        RECT  5.920 2.080 6.200 2.540 ;
        RECT  4.920 1.840 5.120 2.540 ;
        RECT  3.800 2.080 4.080 2.540 ;
        RECT  1.660 2.080 1.940 2.540 ;
        RECT  0.640 1.870 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.160 -0.140 8.360 0.670 ;
        RECT  7.080 -0.140 7.280 0.670 ;
        RECT  5.920 -0.140 6.200 0.500 ;
        RECT  3.980 -0.140 4.140 0.600 ;
        RECT  0.660 -0.140 0.860 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.680 1.600 ;
        RECT  0.140 0.320 0.340 2.010 ;
        RECT  2.360 0.320 3.820 0.480 ;
        RECT  3.660 0.320 3.820 0.920 ;
        RECT  3.660 0.760 4.400 0.920 ;
        RECT  4.200 0.760 4.400 1.600 ;
        RECT  2.840 1.440 4.400 1.600 ;
        RECT  1.220 1.760 3.000 1.920 ;
        RECT  2.840 1.440 3.000 2.050 ;
        RECT  2.640 1.760 3.000 2.050 ;
        RECT  1.220 1.760 1.420 2.080 ;
        RECT  4.580 0.360 5.160 0.560 ;
        RECT  5.740 1.000 5.940 1.540 ;
        RECT  4.580 1.380 5.940 1.540 ;
        RECT  4.580 0.360 4.740 1.920 ;
        RECT  3.360 1.760 4.740 1.920 ;
        RECT  3.360 1.760 3.640 2.080 ;
        RECT  5.400 0.320 5.600 0.820 ;
        RECT  5.400 0.660 6.260 0.820 ;
        RECT  6.100 0.660 6.260 1.920 ;
        RECT  7.280 0.970 7.480 1.920 ;
        RECT  5.400 1.760 7.480 1.920 ;
        RECT  5.400 1.760 5.600 2.080 ;
        LAYER VTPH ;
        RECT  5.600 1.080 7.400 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.080 ;
        RECT  0.000 0.000 5.600 1.140 ;
        RECT  7.400 0.000 8.800 1.140 ;
    END
END LARSM4HM

MACRO LARSM2HM
    CLASS CORE ;
    FOREIGN LARSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.454  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.500 0.760 1.700 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.660 1.700 1.160 ;
        LAYER ME1 ;
        RECT  1.400 0.700 1.880 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.140 1.280 ;
        RECT  2.060 1.080 3.140 1.280 ;
        RECT  2.060 0.940 2.340 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.280 0.390 7.500 2.080 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.480 0.430 6.760 1.600 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.080 3.960 1.280 ;
        RECT  3.300 0.620 3.500 1.280 ;
        RECT  2.040 0.620 3.500 0.780 ;
        RECT  2.040 0.320 2.200 0.780 ;
        RECT  1.040 0.320 2.200 0.480 ;
        RECT  1.040 0.320 1.240 0.960 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.760 5.180 1.160 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.800 1.480 8.000 2.540 ;
        RECT  5.920 2.080 6.200 2.540 ;
        RECT  4.920 1.840 5.120 2.540 ;
        RECT  3.800 2.080 4.080 2.540 ;
        RECT  1.660 2.080 1.940 2.540 ;
        RECT  0.640 1.870 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.800 -0.140 8.000 0.670 ;
        RECT  5.920 -0.140 6.200 0.500 ;
        RECT  3.980 -0.140 4.140 0.600 ;
        RECT  0.660 -0.140 0.860 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.680 1.600 ;
        RECT  0.140 0.320 0.340 2.050 ;
        RECT  2.360 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  3.660 0.760 4.400 0.920 ;
        RECT  4.200 0.760 4.400 1.600 ;
        RECT  2.840 1.440 4.400 1.600 ;
        RECT  1.220 1.760 3.000 1.920 ;
        RECT  2.840 1.440 3.000 2.050 ;
        RECT  2.640 1.760 3.000 2.050 ;
        RECT  1.220 1.760 1.420 2.080 ;
        RECT  4.580 0.360 5.160 0.560 ;
        RECT  5.740 1.000 5.940 1.480 ;
        RECT  4.580 1.320 5.940 1.480 ;
        RECT  4.580 0.360 4.740 1.920 ;
        RECT  3.360 1.760 4.740 1.920 ;
        RECT  3.360 1.760 3.640 2.080 ;
        RECT  5.360 0.350 5.640 0.840 ;
        RECT  5.360 0.660 6.260 0.840 ;
        RECT  6.100 0.660 6.260 1.920 ;
        RECT  6.920 1.000 7.120 1.920 ;
        RECT  5.320 1.760 7.120 1.920 ;
        LAYER VTPH ;
        RECT  5.600 1.080 7.040 2.400 ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.080 ;
        RECT  0.000 0.000 5.600 1.140 ;
        RECT  7.040 0.000 8.400 1.140 ;
    END
END LARSM2HM

MACRO LARSM1HM
    CLASS CORE ;
    FOREIGN LARSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.115  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.580 0.760 1.780 0.960 ;
        LAYER ME2 ;
        RECT  1.580 0.660 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.480 0.700 1.940 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.180 1.280 ;
        RECT  2.980 1.000 3.180 1.280 ;
        RECT  2.140 1.080 3.180 1.280 ;
        RECT  2.140 0.940 2.420 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.040 0.840 7.500 1.160 ;
        RECT  7.040 0.350 7.240 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.272  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.430 6.800 1.600 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.340 1.080 4.020 1.280 ;
        RECT  3.340 0.620 3.500 1.280 ;
        RECT  2.100 0.620 3.500 0.780 ;
        RECT  2.100 0.320 2.300 0.780 ;
        RECT  1.120 0.320 2.300 0.480 ;
        RECT  1.120 0.320 1.320 0.960 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.920 0.840 5.500 1.160 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.560 1.530 7.760 2.540 ;
        RECT  5.960 2.080 6.240 2.540 ;
        RECT  4.960 1.760 5.160 2.540 ;
        RECT  3.820 2.080 4.100 2.540 ;
        RECT  1.740 2.080 2.020 2.540 ;
        RECT  0.720 1.870 1.000 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.560 -0.140 7.760 0.630 ;
        RECT  5.960 -0.140 6.240 0.320 ;
        RECT  4.020 -0.140 4.180 0.600 ;
        RECT  0.740 -0.140 0.940 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.760 1.600 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.460 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  3.660 0.760 4.440 0.920 ;
        RECT  4.280 0.760 4.440 1.600 ;
        RECT  2.920 1.440 4.440 1.600 ;
        RECT  1.300 1.760 3.080 1.920 ;
        RECT  2.920 1.440 3.080 2.070 ;
        RECT  2.680 1.760 3.080 2.070 ;
        RECT  1.300 1.760 1.500 2.080 ;
        RECT  4.600 0.360 5.200 0.560 ;
        RECT  5.780 1.000 5.980 1.480 ;
        RECT  4.600 1.320 5.980 1.480 ;
        RECT  4.600 0.360 4.760 1.920 ;
        RECT  3.460 1.760 4.760 1.920 ;
        RECT  3.460 1.760 3.660 2.100 ;
        RECT  5.400 0.350 5.680 0.660 ;
        RECT  5.400 0.480 6.300 0.660 ;
        RECT  6.140 0.480 6.300 1.920 ;
        RECT  5.360 1.760 6.660 1.920 ;
        RECT  6.500 1.760 6.660 2.100 ;
        RECT  6.500 1.940 7.080 2.100 ;
        LAYER VTPH ;
        RECT  5.640 1.080 7.080 2.400 ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.080 ;
        RECT  0.000 0.000 5.640 1.140 ;
        RECT  7.080 0.000 8.000 1.140 ;
    END
END LARSM1HM

MACRO LARSM0HM
    CLASS CORE ;
    FOREIGN LARSM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.115  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.580 0.760 1.780 0.960 ;
        LAYER ME2 ;
        RECT  1.580 0.660 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.480 0.700 1.940 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.180 1.280 ;
        RECT  2.980 1.000 3.180 1.280 ;
        RECT  2.140 1.080 3.180 1.280 ;
        RECT  2.140 0.940 2.420 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.221  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.080 0.840 7.500 1.160 ;
        RECT  7.080 0.360 7.280 1.720 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.225  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.430 6.840 1.600 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.340 1.080 4.020 1.280 ;
        RECT  3.340 0.620 3.500 1.280 ;
        RECT  2.100 0.620 3.500 0.780 ;
        RECT  2.100 0.320 2.300 0.780 ;
        RECT  1.120 0.320 2.300 0.480 ;
        RECT  1.120 0.320 1.320 0.960 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.920 0.840 5.500 1.160 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.600 1.530 7.800 2.540 ;
        RECT  6.000 2.080 6.280 2.540 ;
        RECT  4.960 1.700 5.160 2.540 ;
        RECT  3.820 2.080 4.100 2.540 ;
        RECT  1.740 2.080 2.020 2.540 ;
        RECT  0.720 1.870 1.000 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.600 -0.140 7.800 0.640 ;
        RECT  6.000 -0.140 6.280 0.320 ;
        RECT  4.020 -0.140 4.180 0.600 ;
        RECT  0.740 -0.140 0.940 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.760 1.600 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.460 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  3.660 0.760 4.440 0.920 ;
        RECT  4.280 0.760 4.440 1.600 ;
        RECT  2.920 1.440 4.440 1.600 ;
        RECT  1.300 1.760 3.080 1.920 ;
        RECT  2.920 1.440 3.080 2.070 ;
        RECT  2.680 1.760 3.080 2.070 ;
        RECT  1.300 1.760 1.500 2.080 ;
        RECT  4.600 0.330 5.200 0.530 ;
        RECT  5.820 1.000 6.020 1.480 ;
        RECT  4.600 1.320 6.020 1.480 ;
        RECT  4.600 0.330 4.760 1.920 ;
        RECT  3.460 1.760 4.760 1.920 ;
        RECT  3.460 1.760 3.660 2.100 ;
        RECT  5.440 0.380 5.640 0.660 ;
        RECT  5.440 0.480 6.340 0.660 ;
        RECT  6.180 0.480 6.340 1.920 ;
        RECT  5.360 1.760 6.700 1.920 ;
        RECT  6.540 1.760 6.700 2.100 ;
        RECT  6.540 1.940 7.120 2.100 ;
        LAYER VTPH ;
        RECT  5.640 1.080 7.120 2.400 ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.080 ;
        RECT  0.000 0.000 5.640 1.140 ;
        RECT  7.120 0.000 8.000 1.140 ;
    END
END LARSM0HM

MACRO LAQRSM4HM
    CLASS CORE ;
    FOREIGN LAQRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.454  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.500 0.760 1.700 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.660 1.700 1.160 ;
        LAYER ME1 ;
        RECT  1.400 0.700 1.880 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.140 1.280 ;
        RECT  2.060 1.080 3.140 1.280 ;
        RECT  2.060 0.960 2.340 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.480 0.430 6.760 2.100 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.080 3.960 1.280 ;
        RECT  3.300 0.640 3.500 1.280 ;
        RECT  2.040 0.640 3.500 0.800 ;
        RECT  2.040 0.320 2.200 0.800 ;
        RECT  1.040 0.320 2.200 0.480 ;
        RECT  1.040 0.320 1.240 0.940 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.760 5.180 1.160 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  7.040 1.450 7.320 2.540 ;
        RECT  5.920 2.080 6.200 2.540 ;
        RECT  4.920 1.840 5.120 2.540 ;
        RECT  3.800 2.080 4.080 2.540 ;
        RECT  1.660 2.080 1.940 2.540 ;
        RECT  0.640 1.870 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.080 -0.140 7.280 0.670 ;
        RECT  5.920 -0.140 6.200 0.500 ;
        RECT  3.980 -0.140 4.140 0.600 ;
        RECT  0.660 -0.140 0.860 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.680 1.600 ;
        RECT  0.140 0.320 0.340 2.010 ;
        RECT  2.360 0.320 3.820 0.480 ;
        RECT  3.660 0.320 3.820 0.920 ;
        RECT  3.660 0.760 4.400 0.920 ;
        RECT  4.200 0.760 4.400 1.600 ;
        RECT  2.840 1.440 4.400 1.600 ;
        RECT  1.220 1.760 3.000 1.920 ;
        RECT  2.840 1.440 3.000 2.050 ;
        RECT  2.640 1.760 3.000 2.050 ;
        RECT  1.220 1.760 1.420 2.080 ;
        RECT  4.580 0.360 5.160 0.560 ;
        RECT  5.580 1.000 5.780 1.540 ;
        RECT  4.580 1.380 5.780 1.540 ;
        RECT  4.580 0.360 4.740 1.920 ;
        RECT  3.360 1.760 4.740 1.920 ;
        RECT  3.360 1.760 3.640 2.080 ;
        RECT  5.400 0.320 5.600 0.820 ;
        RECT  5.400 0.660 6.310 0.820 ;
        RECT  6.100 0.660 6.310 1.920 ;
        RECT  5.400 1.760 6.310 1.920 ;
        RECT  5.400 1.760 5.600 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END LAQRSM4HM

MACRO LAQRSM2HM
    CLASS CORE ;
    FOREIGN LAQRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.454  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.500 0.760 1.700 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.660 1.700 1.160 ;
        LAYER ME1 ;
        RECT  1.400 0.700 1.880 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.140 1.280 ;
        RECT  2.060 1.080 3.140 1.280 ;
        RECT  2.060 0.940 2.340 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.480 0.430 6.760 2.060 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.080 3.960 1.280 ;
        RECT  3.300 0.620 3.500 1.280 ;
        RECT  2.040 0.620 3.500 0.780 ;
        RECT  2.040 0.320 2.200 0.780 ;
        RECT  1.040 0.320 2.200 0.480 ;
        RECT  1.040 0.320 1.240 0.960 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.760 5.180 1.160 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  5.920 2.080 6.200 2.540 ;
        RECT  4.920 1.840 5.120 2.540 ;
        RECT  3.800 2.080 4.080 2.540 ;
        RECT  1.660 2.080 1.940 2.540 ;
        RECT  0.640 1.870 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  5.920 -0.140 6.200 0.500 ;
        RECT  3.980 -0.140 4.140 0.600 ;
        RECT  0.660 -0.140 0.860 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.680 1.600 ;
        RECT  0.140 0.320 0.340 2.050 ;
        RECT  2.360 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  3.660 0.760 4.400 0.920 ;
        RECT  4.200 0.760 4.400 1.600 ;
        RECT  2.840 1.440 4.400 1.600 ;
        RECT  1.220 1.760 3.000 1.920 ;
        RECT  2.840 1.440 3.000 2.050 ;
        RECT  2.640 1.760 3.000 2.050 ;
        RECT  1.220 1.760 1.420 2.080 ;
        RECT  4.580 0.360 5.160 0.560 ;
        RECT  5.420 1.000 5.620 1.480 ;
        RECT  4.580 1.320 5.620 1.480 ;
        RECT  4.580 0.360 4.740 1.920 ;
        RECT  3.360 1.760 4.740 1.920 ;
        RECT  3.360 1.760 3.640 2.080 ;
        RECT  5.360 0.350 5.640 0.840 ;
        RECT  5.360 0.660 6.260 0.840 ;
        RECT  6.100 0.660 6.260 1.920 ;
        RECT  5.320 1.760 6.260 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END LAQRSM2HM

MACRO LAQRSM1HM
    CLASS CORE ;
    FOREIGN LAQRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.115  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.580 0.760 1.780 0.960 ;
        LAYER ME1 ;
        RECT  1.480 0.700 1.940 0.960 ;
        LAYER ME2 ;
        RECT  1.580 0.660 1.900 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.180 1.280 ;
        RECT  2.980 1.000 3.180 1.280 ;
        RECT  2.140 1.080 3.180 1.280 ;
        RECT  2.140 0.940 2.420 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.430 6.800 1.730 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.340 1.080 4.020 1.280 ;
        RECT  3.340 0.620 3.500 1.280 ;
        RECT  2.100 0.620 3.500 0.780 ;
        RECT  2.100 0.320 2.300 0.780 ;
        RECT  1.120 0.320 2.300 0.480 ;
        RECT  1.120 0.320 1.320 0.960 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.240 1.140 5.500 1.560 ;
        RECT  4.920 1.140 5.500 1.480 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  5.960 2.080 6.240 2.540 ;
        RECT  4.960 1.760 5.160 2.540 ;
        RECT  3.820 2.080 4.100 2.540 ;
        RECT  1.740 2.080 2.020 2.540 ;
        RECT  0.720 1.870 1.000 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  5.960 -0.140 6.240 0.320 ;
        RECT  4.020 -0.140 4.180 0.600 ;
        RECT  0.740 -0.140 0.940 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.760 1.600 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.460 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  3.660 0.760 4.440 0.920 ;
        RECT  4.280 0.760 4.440 1.600 ;
        RECT  2.920 1.440 4.440 1.600 ;
        RECT  1.300 1.760 3.080 1.920 ;
        RECT  2.920 1.440 3.080 2.070 ;
        RECT  2.680 1.760 3.080 2.070 ;
        RECT  1.300 1.760 1.500 2.080 ;
        RECT  4.600 0.360 5.200 0.560 ;
        RECT  4.600 0.800 5.620 0.960 ;
        RECT  4.600 0.360 4.760 1.920 ;
        RECT  3.460 1.760 4.760 1.920 ;
        RECT  3.460 1.760 3.660 2.100 ;
        RECT  5.400 0.350 5.680 0.640 ;
        RECT  5.400 0.480 6.300 0.640 ;
        RECT  6.140 0.480 6.300 1.920 ;
        RECT  5.360 1.760 6.300 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END LAQRSM1HM

MACRO LAQRSM0HM
    CLASS CORE ;
    FOREIGN LAQRSM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.115  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.580 0.760 1.780 0.960 ;
        LAYER ME2 ;
        RECT  1.580 0.660 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.480 0.700 1.940 0.960 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.120 3.180 1.280 ;
        RECT  2.980 1.000 3.180 1.280 ;
        RECT  2.140 1.080 3.180 1.280 ;
        RECT  2.140 0.940 2.420 1.280 ;
        RECT  0.500 0.840 0.700 1.280 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.460 0.430 6.800 1.850 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.340 1.080 4.020 1.280 ;
        RECT  3.340 0.620 3.500 1.280 ;
        RECT  2.100 0.620 3.500 0.780 ;
        RECT  2.100 0.320 2.300 0.780 ;
        RECT  1.120 0.320 2.300 0.480 ;
        RECT  1.120 0.320 1.320 0.960 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.240 1.200 5.500 1.560 ;
        RECT  4.920 1.200 5.500 1.540 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.000 1.610 6.220 2.540 ;
        RECT  4.960 1.700 5.160 2.540 ;
        RECT  3.840 2.080 4.120 2.540 ;
        RECT  1.740 2.080 2.020 2.540 ;
        RECT  0.720 1.870 1.000 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.020 -0.140 6.240 0.670 ;
        RECT  4.020 -0.140 4.180 0.600 ;
        RECT  0.740 -0.140 0.940 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 2.760 1.600 ;
        RECT  0.140 0.320 0.340 2.080 ;
        RECT  2.460 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  3.660 0.760 4.440 0.920 ;
        RECT  4.280 0.760 4.440 1.600 ;
        RECT  2.920 1.440 4.440 1.600 ;
        RECT  1.300 1.760 3.080 1.920 ;
        RECT  2.920 1.440 3.080 2.070 ;
        RECT  2.680 1.760 3.080 2.070 ;
        RECT  1.300 1.760 1.500 2.080 ;
        RECT  4.600 0.330 5.090 0.530 ;
        RECT  4.600 0.800 5.390 0.960 ;
        RECT  4.600 0.330 4.760 1.920 ;
        RECT  3.420 1.760 4.760 1.920 ;
        RECT  3.420 1.760 3.680 2.100 ;
        RECT  5.330 0.300 5.530 0.640 ;
        RECT  5.330 0.460 5.830 0.640 ;
        RECT  5.670 1.000 6.210 1.280 ;
        RECT  5.670 0.460 5.830 1.920 ;
        RECT  5.360 1.760 5.830 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END LAQRSM0HM

MACRO LAQM4HM
    CLASS CORE ;
    FOREIGN LAQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.720 2.160 1.100 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.502  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.060 0.840 5.500 1.160 ;
        RECT  5.060 0.840 5.340 2.100 ;
        RECT  5.060 0.340 5.280 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.640 1.370 5.840 2.540 ;
        RECT  4.520 1.940 4.720 2.540 ;
        RECT  3.510 1.880 3.720 2.540 ;
        RECT  1.700 1.580 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.640 -0.140 5.810 0.760 ;
        RECT  4.570 -0.140 4.770 0.670 ;
        RECT  3.550 -0.140 3.750 0.580 ;
        RECT  1.720 -0.140 1.920 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.320 0.660 2.640 0.940 ;
        RECT  1.280 1.260 2.480 1.420 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.320 0.660 2.480 2.030 ;
        RECT  2.320 1.870 3.320 2.030 ;
        RECT  2.500 0.340 3.060 0.500 ;
        RECT  2.900 0.340 3.060 1.290 ;
        RECT  2.740 1.070 4.110 1.290 ;
        RECT  2.740 1.070 2.900 1.710 ;
        RECT  4.100 0.380 4.260 0.910 ;
        RECT  3.240 0.750 4.430 0.910 ;
        RECT  4.270 0.750 4.430 1.680 ;
        RECT  4.040 1.520 4.430 1.680 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.260 2.400 ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.260 0.000 6.000 1.140 ;
    END
END LAQM4HM

MACRO LAQM2HM
    CLASS CORE ;
    FOREIGN LAQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.750 0.900 5.250 1.100 ;
        RECT  4.750 0.900 4.990 2.100 ;
        RECT  4.750 0.380 4.910 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.270 1.380 5.430 2.540 ;
        RECT  3.700 1.500 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.250 -0.140 5.450 0.700 ;
        RECT  3.540 -0.140 3.740 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.100 ;
        RECT  2.460 1.940 3.280 2.100 ;
        RECT  2.540 0.340 3.080 0.500 ;
        RECT  2.920 0.340 3.080 1.230 ;
        RECT  2.780 1.070 4.260 1.230 ;
        RECT  2.780 1.070 2.940 1.740 ;
        RECT  4.020 0.340 4.300 0.910 ;
        RECT  3.240 0.750 4.580 0.910 ;
        RECT  4.420 0.750 4.580 1.710 ;
        RECT  4.140 1.550 4.580 1.710 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 5.600 1.140 ;
    END
END LAQM2HM

MACRO LAQM1HM
    CLASS CORE ;
    FOREIGN LAQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.760 0.900 5.260 1.100 ;
        RECT  4.760 0.470 4.920 1.780 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.280 1.640 5.480 2.540 ;
        RECT  3.700 1.500 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.260 -0.140 5.460 0.740 ;
        RECT  3.540 -0.140 3.740 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.100 ;
        RECT  2.460 1.940 3.280 2.100 ;
        RECT  2.540 0.340 3.080 0.500 ;
        RECT  2.920 0.340 3.080 1.230 ;
        RECT  2.780 1.070 4.270 1.230 ;
        RECT  2.780 1.070 2.940 1.740 ;
        RECT  4.020 0.340 4.300 0.910 ;
        RECT  3.240 0.750 4.590 0.910 ;
        RECT  4.430 0.750 4.590 1.710 ;
        RECT  4.140 1.550 4.590 1.710 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 5.600 1.140 ;
    END
END LAQM1HM

MACRO LAQM0HM
    CLASS CORE ;
    FOREIGN LAQM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.245  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.720 0.900 5.260 1.100 ;
        RECT  4.720 0.460 4.920 1.780 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.280 1.640 5.480 2.540 ;
        RECT  3.700 1.500 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.260 -0.140 5.460 0.740 ;
        RECT  3.540 -0.140 3.740 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.100 ;
        RECT  2.460 1.940 3.280 2.100 ;
        RECT  2.540 0.340 3.080 0.500 ;
        RECT  2.920 0.340 3.080 1.230 ;
        RECT  2.780 1.070 4.230 1.230 ;
        RECT  2.780 1.070 2.940 1.740 ;
        RECT  4.020 0.340 4.300 0.910 ;
        RECT  3.240 0.750 4.550 0.910 ;
        RECT  4.390 0.750 4.550 1.710 ;
        RECT  4.140 1.550 4.550 1.710 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 5.600 1.140 ;
    END
END LAQM0HM

MACRO LAM4HM
    CLASS CORE ;
    FOREIGN LAM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.550  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.200 0.420 5.500 0.760 ;
        RECT  5.200 0.420 5.360 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.670 6.700 1.600 ;
        RECT  6.340 1.400 6.540 2.100 ;
        RECT  6.260 0.670 6.700 0.870 ;
        RECT  6.260 0.420 6.460 0.870 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.860 1.760 7.060 2.540 ;
        RECT  5.840 1.720 6.040 2.540 ;
        RECT  4.520 1.940 4.720 2.540 ;
        RECT  3.640 1.880 3.850 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.740 -0.140 7.020 0.510 ;
        RECT  5.740 -0.140 5.940 0.700 ;
        RECT  4.700 -0.140 4.900 0.590 ;
        RECT  3.700 -0.140 3.900 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.030 ;
        RECT  2.460 1.870 3.360 2.030 ;
        RECT  2.540 0.340 3.100 0.500 ;
        RECT  2.940 0.340 3.100 1.230 ;
        RECT  2.780 1.070 4.300 1.230 ;
        RECT  2.780 1.070 2.940 1.710 ;
        RECT  4.240 0.380 4.400 0.910 ;
        RECT  3.280 0.750 4.660 0.910 ;
        RECT  5.800 1.040 6.340 1.240 ;
        RECT  4.500 0.750 4.660 1.680 ;
        RECT  5.800 1.040 5.960 1.560 ;
        RECT  5.520 1.400 5.960 1.560 ;
        RECT  4.120 1.520 5.040 1.680 ;
        RECT  4.880 1.520 5.040 2.100 ;
        RECT  5.520 1.400 5.680 2.100 ;
        RECT  4.880 1.940 5.680 2.100 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 7.200 1.140 ;
    END
END LAM4HM

MACRO LAM2HM
    CLASS CORE ;
    FOREIGN LAM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.770 0.900 5.270 1.100 ;
        RECT  4.770 0.380 4.930 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.930 0.440 6.130 2.100 ;
        RECT  5.700 0.440 6.130 0.760 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.410 1.640 5.570 2.540 ;
        RECT  3.700 1.500 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.270 -0.140 5.470 0.700 ;
        RECT  3.540 -0.140 3.740 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.100 ;
        RECT  2.460 1.940 3.280 2.100 ;
        RECT  2.540 0.340 3.080 0.500 ;
        RECT  2.920 0.340 3.080 1.230 ;
        RECT  2.780 1.070 4.280 1.230 ;
        RECT  2.780 1.070 2.940 1.740 ;
        RECT  4.020 0.340 4.300 0.910 ;
        RECT  3.240 0.750 4.600 0.910 ;
        RECT  5.590 0.960 5.750 1.480 ;
        RECT  5.090 1.320 5.750 1.480 ;
        RECT  4.140 1.550 4.600 1.710 ;
        RECT  4.440 0.750 4.600 2.100 ;
        RECT  5.090 1.320 5.250 2.100 ;
        RECT  4.440 1.940 5.250 2.100 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 6.400 1.140 ;
    END
END LAM2HM

MACRO LAM1HM
    CLASS CORE ;
    FOREIGN LAM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.770 0.900 5.270 1.100 ;
        RECT  4.770 0.470 4.930 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.930 0.440 6.130 1.820 ;
        RECT  5.700 0.440 6.130 0.760 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.410 1.640 5.610 2.540 ;
        RECT  3.700 1.500 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.270 -0.140 5.470 0.740 ;
        RECT  3.540 -0.140 3.740 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.100 ;
        RECT  2.460 1.940 3.280 2.100 ;
        RECT  2.540 0.340 3.080 0.500 ;
        RECT  2.920 0.340 3.080 1.230 ;
        RECT  2.780 1.070 4.280 1.230 ;
        RECT  2.780 1.070 2.940 1.740 ;
        RECT  4.020 0.340 4.300 0.910 ;
        RECT  3.240 0.750 4.600 0.910 ;
        RECT  5.590 0.960 5.750 1.480 ;
        RECT  5.090 1.320 5.750 1.480 ;
        RECT  4.140 1.550 4.600 1.710 ;
        RECT  4.440 0.750 4.600 2.100 ;
        RECT  5.090 1.320 5.250 2.100 ;
        RECT  4.440 1.940 5.250 2.100 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 6.400 1.140 ;
    END
END LAM1HM

MACRO LAM0HM
    CLASS CORE ;
    FOREIGN LAM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.245  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.730 0.900 5.270 1.100 ;
        RECT  4.730 0.460 4.930 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.245  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.930 0.440 6.130 1.850 ;
        RECT  5.700 0.440 6.130 0.760 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.410 1.640 5.610 2.540 ;
        RECT  3.700 1.500 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.270 -0.140 5.470 0.740 ;
        RECT  3.540 -0.140 3.740 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  2.460 0.660 2.680 0.940 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 0.660 2.620 2.100 ;
        RECT  2.460 1.940 3.280 2.100 ;
        RECT  2.540 0.340 3.080 0.500 ;
        RECT  2.920 0.340 3.080 1.230 ;
        RECT  2.780 1.070 4.240 1.230 ;
        RECT  2.780 1.070 2.940 1.740 ;
        RECT  4.020 0.340 4.300 0.910 ;
        RECT  3.240 0.750 4.560 0.910 ;
        RECT  5.590 0.960 5.750 1.480 ;
        RECT  5.090 1.320 5.750 1.480 ;
        RECT  4.140 1.550 4.560 1.710 ;
        RECT  4.400 0.750 4.560 2.100 ;
        RECT  5.090 1.320 5.250 2.100 ;
        RECT  4.400 1.940 5.250 2.100 ;
        LAYER VTPH ;
        RECT  1.400 1.060 3.300 2.400 ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.060 ;
        RECT  0.000 0.000 1.400 1.140 ;
        RECT  3.300 0.000 6.400 1.140 ;
    END
END LAM0HM

MACRO LAGCESM8HM
    CLASS CORE ;
    FOREIGN LAGCESM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.223  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.700 1.040 6.120 1.240 ;
        RECT  5.700 0.840 5.900 1.240 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.825  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.580 0.660 8.820 0.860 ;
        RECT  8.620 0.310 8.820 0.860 ;
        RECT  8.100 0.660 8.300 2.100 ;
        RECT  7.060 1.420 8.300 1.620 ;
        RECT  7.580 0.310 7.780 0.860 ;
        RECT  7.060 1.420 7.260 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.620 1.800 8.820 2.540 ;
        RECT  7.580 1.800 7.780 2.540 ;
        RECT  6.540 1.780 6.740 2.540 ;
        RECT  5.500 1.720 5.700 2.540 ;
        RECT  4.280 1.630 4.480 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.060 -0.140 8.340 0.500 ;
        RECT  7.060 -0.140 7.260 0.610 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.540 0.840 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.820 0.980 4.980 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.300 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  6.140 0.300 6.300 0.880 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.140 0.720 6.540 0.880 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  6.380 0.720 6.540 1.260 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.460 0.400 6.860 0.560 ;
        RECT  6.700 1.020 7.880 1.180 ;
        RECT  6.700 0.400 6.860 1.620 ;
        RECT  6.180 1.460 6.860 1.620 ;
        RECT  6.180 1.460 6.380 1.920 ;
        RECT  5.980 1.720 6.380 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.200 1.140 ;
    END
END LAGCESM8HM

MACRO LAGCESM6HM
    CLASS CORE ;
    FOREIGN LAGCESM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.223  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.700 1.040 6.120 1.240 ;
        RECT  5.700 0.840 5.900 1.240 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.675  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.080 1.420 8.300 2.100 ;
        RECT  8.100 0.660 8.300 2.100 ;
        RECT  7.540 0.660 8.300 0.860 ;
        RECT  7.020 1.420 8.300 1.620 ;
        RECT  7.540 0.360 7.740 0.860 ;
        RECT  7.020 1.420 7.220 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.540 1.800 7.740 2.540 ;
        RECT  6.500 1.780 6.700 2.540 ;
        RECT  5.460 1.720 5.660 2.540 ;
        RECT  4.280 1.630 4.480 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  8.020 -0.140 8.300 0.500 ;
        RECT  7.020 -0.140 7.220 0.630 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.540 0.840 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.820 0.980 4.980 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.300 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  6.140 0.300 6.300 0.880 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.140 0.720 6.540 0.880 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  6.380 0.720 6.540 1.290 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.460 0.400 6.860 0.560 ;
        RECT  6.700 1.020 7.840 1.180 ;
        RECT  6.700 0.400 6.860 1.620 ;
        RECT  6.140 1.460 6.860 1.620 ;
        RECT  6.140 1.460 6.340 1.920 ;
        RECT  5.940 1.720 6.340 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END LAGCESM6HM

MACRO LAGCESM4HM
    CLASS CORE ;
    FOREIGN LAGCESM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.223  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.700 1.040 6.120 1.240 ;
        RECT  5.700 0.840 5.900 1.240 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.020 1.420 7.900 1.620 ;
        RECT  7.700 0.460 7.900 1.620 ;
        RECT  7.500 0.460 7.900 0.660 ;
        RECT  7.020 1.420 7.220 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.540 1.800 7.740 2.540 ;
        RECT  6.500 1.780 6.700 2.540 ;
        RECT  5.460 1.720 5.660 2.540 ;
        RECT  4.280 1.630 4.480 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.020 -0.140 7.220 0.700 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.540 0.840 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.820 0.980 4.980 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.300 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  6.140 0.300 6.300 0.880 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.140 0.720 6.540 0.880 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  6.380 0.720 6.540 1.290 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.460 0.400 6.860 0.560 ;
        RECT  6.700 1.020 7.480 1.180 ;
        RECT  6.700 0.400 6.860 1.620 ;
        RECT  6.140 1.460 6.860 1.620 ;
        RECT  6.140 1.460 6.340 1.920 ;
        RECT  5.940 1.720 6.340 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END LAGCESM4HM

MACRO LAGCESM3HM
    CLASS CORE ;
    FOREIGN LAGCESM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.223  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.700 1.040 6.120 1.240 ;
        RECT  5.700 0.840 5.900 1.240 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.350  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.020 1.420 7.900 1.620 ;
        RECT  7.700 0.530 7.900 1.620 ;
        RECT  7.500 0.530 7.900 0.730 ;
        RECT  7.020 1.420 7.220 2.000 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.540 1.800 7.740 2.540 ;
        RECT  6.500 1.780 6.700 2.540 ;
        RECT  5.460 1.720 5.660 2.540 ;
        RECT  4.280 1.630 4.480 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.020 -0.140 7.220 0.760 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.540 0.840 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.820 0.980 4.980 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.300 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  6.140 0.300 6.300 0.880 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.140 0.720 6.540 0.880 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  6.380 0.720 6.540 1.290 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.460 0.400 6.860 0.560 ;
        RECT  6.700 1.100 7.480 1.260 ;
        RECT  6.700 0.400 6.860 1.620 ;
        RECT  6.140 1.460 6.860 1.620 ;
        RECT  6.140 1.460 6.340 1.920 ;
        RECT  5.940 1.720 6.340 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END LAGCESM3HM

MACRO LAGCESM2HM
    CLASS CORE ;
    FOREIGN LAGCESM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.070 1.220 6.240 1.420 ;
        RECT  5.300 1.220 5.500 1.560 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.326  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.880 0.440 7.100 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.300 1.900 6.580 2.540 ;
        RECT  5.300 1.790 5.500 2.540 ;
        RECT  4.300 1.630 4.500 2.540 ;
        RECT  2.460 1.860 2.740 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.300 -0.140 6.580 0.660 ;
        RECT  2.880 -0.140 3.080 0.380 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.720 0.460 ;
        RECT  2.560 0.300 2.720 0.700 ;
        RECT  2.560 0.540 3.060 0.700 ;
        RECT  2.900 0.540 3.060 1.060 ;
        RECT  2.900 0.900 3.320 1.060 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.590 1.500 1.900 1.780 ;
        RECT  3.800 0.620 4.180 0.820 ;
        RECT  2.060 0.640 2.400 0.860 ;
        RECT  1.270 1.060 1.540 1.340 ;
        RECT  2.060 1.540 3.060 1.700 ;
        RECT  2.900 1.540 3.060 2.040 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  3.800 0.620 3.960 2.040 ;
        RECT  2.900 1.880 3.960 2.040 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  4.750 0.690 5.220 0.850 ;
        RECT  4.140 0.980 4.910 1.140 ;
        RECT  4.140 0.980 4.300 1.410 ;
        RECT  4.750 0.690 4.910 1.850 ;
        RECT  4.750 1.690 5.100 1.850 ;
        RECT  3.480 0.300 5.360 0.460 ;
        RECT  2.460 1.060 2.660 1.380 ;
        RECT  3.480 0.300 3.640 1.380 ;
        RECT  2.460 1.220 3.640 1.380 ;
        RECT  3.220 1.220 3.420 1.720 ;
        RECT  5.520 0.430 5.680 1.000 ;
        RECT  5.520 0.840 6.700 1.000 ;
        RECT  6.540 0.840 6.700 1.740 ;
        RECT  5.840 1.580 6.700 1.740 ;
        RECT  5.840 1.580 6.000 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.160 2.400 ;
        RECT  5.480 1.140 7.200 2.400 ;
        RECT  0.000 1.220 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
        RECT  4.160 0.000 5.480 1.220 ;
    END
END LAGCESM2HM

MACRO LAGCESM20HM
    CLASS CORE ;
    FOREIGN LAGCESM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.425  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.640 1.230 7.820 1.390 ;
        RECT  5.640 0.840 5.900 1.390 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.039  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.080 1.410 13.280 2.100 ;
        RECT  8.920 1.420 13.280 1.620 ;
        RECT  10.850 1.410 13.280 1.620 ;
        RECT  9.440 0.660 12.760 0.860 ;
        RECT  12.560 0.320 12.760 0.860 ;
        RECT  12.040 1.410 12.240 2.050 ;
        RECT  11.520 0.320 11.720 0.860 ;
        RECT  11.000 1.410 11.200 2.050 ;
        RECT  10.850 0.660 11.150 1.620 ;
        RECT  10.480 0.320 10.680 0.860 ;
        RECT  9.960 1.420 10.160 2.050 ;
        RECT  9.440 0.320 9.640 0.860 ;
        RECT  8.920 1.420 9.120 2.060 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.560 1.800 12.760 2.540 ;
        RECT  11.520 1.800 11.720 2.540 ;
        RECT  10.480 1.800 10.680 2.540 ;
        RECT  9.440 1.800 9.640 2.540 ;
        RECT  8.360 1.870 8.640 2.540 ;
        RECT  7.320 1.870 7.600 2.540 ;
        RECT  6.280 1.870 6.560 2.540 ;
        RECT  5.280 1.800 5.480 2.540 ;
        RECT  4.280 1.630 4.480 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  13.080 -0.140 13.280 0.570 ;
        RECT  12.000 -0.140 12.280 0.500 ;
        RECT  10.960 -0.140 11.240 0.500 ;
        RECT  9.920 -0.140 10.200 0.500 ;
        RECT  8.920 -0.140 9.120 0.600 ;
        RECT  7.360 -0.140 7.640 0.430 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.820 0.980 4.980 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.320 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.160 0.300 6.320 1.070 ;
        RECT  6.160 0.910 8.280 1.070 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  8.120 0.910 8.280 1.320 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.540 0.400 6.700 0.750 ;
        RECT  8.300 0.340 8.460 0.750 ;
        RECT  6.540 0.590 8.600 0.750 ;
        RECT  8.440 1.020 10.600 1.180 ;
        RECT  8.440 0.590 8.600 1.710 ;
        RECT  5.800 1.550 8.600 1.710 ;
        RECT  5.800 1.550 6.000 1.970 ;
        RECT  6.840 1.550 7.040 1.970 ;
        RECT  7.880 1.550 8.080 1.970 ;
        RECT  11.400 1.020 12.840 1.180 ;
        LAYER VTPH ;
        RECT  8.000 1.050 12.960 2.400 ;
        RECT  0.000 1.140 4.900 2.400 ;
        RECT  8.000 1.140 13.600 2.400 ;
        RECT  0.000 1.240 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.050 ;
        RECT  0.000 0.000 8.000 1.140 ;
        RECT  12.960 0.000 13.600 1.140 ;
        RECT  4.900 0.000 8.000 1.240 ;
    END
END LAGCESM20HM

MACRO LAGCESM16HM
    CLASS CORE ;
    FOREIGN LAGCESM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.356  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.700 1.200 7.340 1.360 ;
        RECT  7.180 0.900 7.340 1.360 ;
        RECT  5.700 0.840 5.900 1.360 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.647  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.160 1.410 11.360 2.100 ;
        RECT  8.040 1.420 11.360 1.620 ;
        RECT  9.250 1.410 11.360 1.620 ;
        RECT  8.560 0.660 10.840 0.840 ;
        RECT  10.640 0.330 10.840 0.840 ;
        RECT  10.120 1.410 10.320 2.050 ;
        RECT  9.600 0.330 9.800 0.840 ;
        RECT  9.250 0.660 9.550 1.620 ;
        RECT  9.080 1.420 9.280 2.050 ;
        RECT  8.560 0.330 8.760 0.840 ;
        RECT  8.040 1.420 8.240 2.060 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.640 1.800 10.840 2.540 ;
        RECT  9.600 1.800 9.800 2.540 ;
        RECT  8.560 1.800 8.760 2.540 ;
        RECT  7.480 1.840 7.760 2.540 ;
        RECT  6.440 1.840 6.720 2.540 ;
        RECT  5.440 1.800 5.640 2.540 ;
        RECT  4.280 1.630 4.480 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.160 -0.140 11.360 0.600 ;
        RECT  10.080 -0.140 10.360 0.500 ;
        RECT  9.040 -0.140 9.320 0.500 ;
        RECT  8.040 -0.140 8.240 0.610 ;
        RECT  7.320 -0.140 7.600 0.400 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.820 0.980 4.980 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.310 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.150 0.300 6.310 1.040 ;
        RECT  6.150 0.880 6.940 1.040 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.500 0.300 6.660 0.720 ;
        RECT  6.500 0.560 7.720 0.720 ;
        RECT  7.560 1.000 9.000 1.160 ;
        RECT  7.560 0.560 7.720 1.680 ;
        RECT  6.080 1.520 7.720 1.680 ;
        RECT  6.080 1.520 6.280 2.000 ;
        RECT  5.920 1.800 6.280 2.000 ;
        RECT  7.000 1.520 7.200 2.100 ;
        RECT  9.800 1.000 10.880 1.160 ;
        LAYER VTPH ;
        RECT  5.770 1.020 11.040 2.400 ;
        RECT  0.000 1.140 4.260 2.400 ;
        RECT  5.770 1.140 11.600 2.400 ;
        RECT  0.000 1.240 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.020 ;
        RECT  0.000 0.000 5.770 1.140 ;
        RECT  11.040 0.000 11.600 1.140 ;
        RECT  4.260 0.000 5.770 1.240 ;
    END
END LAGCESM16HM

MACRO LAGCESM12HM
    CLASS CORE ;
    FOREIGN LAGCESM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.580 1.200 7.340 1.360 ;
        RECT  7.180 0.900 7.340 1.360 ;
        RECT  5.580 1.140 5.900 1.360 ;
        RECT  5.700 0.840 5.900 1.360 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.204  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.380 0.660 10.660 0.860 ;
        RECT  10.460 0.310 10.660 0.860 ;
        RECT  9.940 1.410 10.140 2.100 ;
        RECT  7.860 1.420 10.140 1.620 ;
        RECT  8.850 1.410 10.140 1.620 ;
        RECT  9.420 0.310 9.620 0.860 ;
        RECT  8.850 0.660 9.150 1.620 ;
        RECT  8.900 0.660 9.100 2.100 ;
        RECT  8.380 0.310 8.580 0.860 ;
        RECT  7.860 1.420 8.060 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 1.110 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  10.460 1.800 10.660 2.540 ;
        RECT  9.420 1.800 9.620 2.540 ;
        RECT  8.380 1.800 8.580 2.540 ;
        RECT  7.300 1.840 7.580 2.540 ;
        RECT  6.260 1.840 6.540 2.540 ;
        RECT  5.260 1.730 5.460 2.540 ;
        RECT  4.260 1.630 4.460 2.540 ;
        RECT  2.460 1.830 2.740 2.540 ;
        RECT  0.260 1.720 0.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  9.900 -0.140 10.180 0.500 ;
        RECT  8.860 -0.140 9.140 0.500 ;
        RECT  7.860 -0.140 8.060 0.610 ;
        RECT  7.340 -0.140 7.620 0.400 ;
        RECT  4.620 -0.140 4.780 0.500 ;
        RECT  2.920 -0.140 3.120 0.560 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.740 0.300 2.760 0.460 ;
        RECT  2.600 0.300 2.760 0.880 ;
        RECT  2.600 0.720 3.200 0.880 ;
        RECT  3.000 0.720 3.200 1.030 ;
        RECT  1.740 0.300 1.900 1.780 ;
        RECT  1.600 1.500 1.900 1.780 ;
        RECT  3.780 0.620 4.140 0.820 ;
        RECT  2.060 0.640 2.440 0.840 ;
        RECT  1.270 1.060 1.580 1.340 ;
        RECT  2.060 1.510 3.060 1.670 ;
        RECT  1.270 1.060 1.430 2.100 ;
        RECT  2.900 1.510 3.060 2.100 ;
        RECT  3.700 1.610 3.940 2.100 ;
        RECT  2.060 0.640 2.220 2.100 ;
        RECT  1.270 1.940 2.220 2.100 ;
        RECT  3.780 0.620 3.940 2.100 ;
        RECT  2.900 1.940 3.940 2.100 ;
        RECT  5.260 0.620 5.420 1.140 ;
        RECT  4.120 0.980 5.420 1.140 ;
        RECT  4.120 0.980 4.280 1.410 ;
        RECT  4.800 0.980 4.960 1.950 ;
        RECT  3.440 0.300 4.460 0.460 ;
        RECT  4.940 0.300 6.360 0.460 ;
        RECT  4.300 0.300 4.460 0.820 ;
        RECT  4.940 0.300 5.100 0.820 ;
        RECT  4.300 0.660 5.100 0.820 ;
        RECT  6.200 0.300 6.360 1.040 ;
        RECT  6.200 0.880 6.960 1.040 ;
        RECT  2.430 1.060 2.630 1.350 ;
        RECT  3.440 0.300 3.600 1.350 ;
        RECT  2.430 1.190 3.600 1.350 ;
        RECT  3.220 1.190 3.420 1.760 ;
        RECT  6.520 0.320 6.720 0.720 ;
        RECT  6.520 0.560 7.660 0.720 ;
        RECT  7.500 1.020 8.680 1.180 ;
        RECT  7.500 0.560 7.660 1.680 ;
        RECT  5.900 1.520 7.660 1.680 ;
        RECT  5.900 1.520 6.100 2.000 ;
        RECT  5.740 1.800 6.100 2.000 ;
        RECT  6.820 1.520 7.020 2.000 ;
        RECT  9.320 1.020 10.400 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.260 2.400 ;
        RECT  5.770 1.140 10.800 2.400 ;
        RECT  0.000 1.240 10.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.800 1.140 ;
        RECT  4.260 0.000 5.770 1.240 ;
    END
END LAGCESM12HM

MACRO LAGCEM8HM
    CLASS CORE ;
    FOREIGN LAGCEM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.266  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 1.080 1.340 ;
        RECT  0.100 0.840 0.300 1.340 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.281  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.410 2.360 0.930 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.560 1.520 11.480 1.680 ;
        RECT  11.320 0.480 11.480 1.680 ;
        RECT  7.960 0.480 11.480 0.640 ;
        RECT  10.320 1.520 10.700 2.060 ;
        RECT  10.460 0.320 10.660 0.640 ;
        RECT  9.160 0.320 9.360 0.640 ;
        RECT  8.560 1.520 8.760 2.020 ;
        RECT  7.960 0.320 8.160 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.120 1.880 11.400 2.540 ;
        RECT  9.440 1.840 9.640 2.540 ;
        RECT  7.380 1.820 7.580 2.540 ;
        RECT  6.180 2.080 6.460 2.540 ;
        RECT  2.980 2.080 3.260 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.160 -0.140 11.440 0.320 ;
        RECT  9.720 -0.140 10.000 0.320 ;
        RECT  8.520 -0.140 8.800 0.320 ;
        RECT  7.380 -0.140 7.540 0.640 ;
        RECT  6.170 -0.140 6.370 0.610 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  1.140 -0.140 1.420 0.550 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.340 1.440 3.910 1.600 ;
        RECT  2.540 0.440 2.740 0.900 ;
        RECT  3.580 0.370 3.780 0.900 ;
        RECT  4.600 0.620 4.920 0.900 ;
        RECT  2.540 0.700 4.920 0.900 ;
        RECT  1.740 1.090 5.020 1.250 ;
        RECT  1.740 0.300 1.940 1.260 ;
        RECT  4.750 1.090 5.020 1.290 ;
        RECT  1.860 1.090 2.060 1.780 ;
        RECT  4.060 0.300 5.340 0.460 ;
        RECT  4.060 0.300 4.340 0.540 ;
        RECT  5.180 0.300 5.340 1.780 ;
        RECT  5.180 0.900 6.510 1.100 ;
        RECT  5.180 0.900 5.360 1.780 ;
        RECT  4.100 1.560 5.360 1.780 ;
        RECT  6.670 0.480 6.870 1.600 ;
        RECT  5.910 1.380 6.870 1.600 ;
        RECT  7.060 0.800 10.780 0.960 ;
        RECT  7.060 0.800 7.260 1.180 ;
        RECT  0.660 0.370 0.860 0.870 ;
        RECT  0.660 0.710 1.500 0.870 ;
        RECT  10.960 0.950 11.160 1.340 ;
        RECT  7.460 1.120 11.160 1.340 ;
        RECT  1.340 0.710 1.500 1.680 ;
        RECT  7.460 1.120 7.620 1.580 ;
        RECT  7.040 1.420 7.620 1.580 ;
        RECT  0.660 1.520 1.700 1.680 ;
        RECT  2.220 1.760 3.580 1.920 ;
        RECT  7.040 1.420 7.200 1.920 ;
        RECT  5.810 1.760 7.200 1.920 ;
        RECT  1.540 1.520 1.700 2.100 ;
        RECT  3.420 1.760 3.580 2.100 ;
        RECT  0.660 1.520 0.860 2.070 ;
        RECT  2.220 1.760 2.380 2.100 ;
        RECT  1.540 1.940 2.380 2.100 ;
        RECT  5.810 1.760 5.970 2.100 ;
        RECT  3.420 1.940 5.970 2.100 ;
        LAYER VTPH ;
        RECT  2.200 1.080 4.040 2.400 ;
        RECT  6.320 1.060 7.290 2.400 ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.060 ;
        RECT  0.000 0.000 6.320 1.080 ;
        RECT  0.000 0.000 2.200 1.140 ;
        RECT  4.040 0.000 6.320 1.140 ;
        RECT  7.290 0.000 11.600 1.140 ;
    END
END LAGCEM8HM

MACRO LAGCEM6HM
    CLASS CORE ;
    FOREIGN LAGCEM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.199  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 1.080 1.340 ;
        RECT  0.100 0.840 0.300 1.340 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.226  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.410 2.360 0.930 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.740  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.920 1.520 10.300 2.060 ;
        RECT  10.080 0.480 10.300 2.060 ;
        RECT  7.960 0.480 10.300 0.640 ;
        RECT  8.240 1.520 10.300 1.680 ;
        RECT  9.040 0.320 9.240 0.640 ;
        RECT  8.240 1.520 8.440 2.020 ;
        RECT  7.960 0.320 8.160 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.080 1.840 9.280 2.540 ;
        RECT  7.380 1.820 7.580 2.540 ;
        RECT  6.180 2.080 6.460 2.540 ;
        RECT  2.980 2.080 3.260 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.790 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.600 -0.140 9.880 0.320 ;
        RECT  8.480 -0.140 8.760 0.320 ;
        RECT  7.380 -0.140 7.540 0.640 ;
        RECT  6.170 -0.140 6.370 0.610 ;
        RECT  3.020 -0.140 3.300 0.540 ;
        RECT  1.140 -0.140 1.420 0.530 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.340 1.440 3.910 1.600 ;
        RECT  2.540 0.440 2.740 0.900 ;
        RECT  3.580 0.370 3.780 0.900 ;
        RECT  4.600 0.620 4.920 0.900 ;
        RECT  2.540 0.700 4.920 0.900 ;
        RECT  1.740 1.090 5.020 1.250 ;
        RECT  4.750 1.090 5.020 1.290 ;
        RECT  1.740 0.300 1.940 1.350 ;
        RECT  1.860 1.090 2.060 1.780 ;
        RECT  4.060 0.300 5.340 0.460 ;
        RECT  4.060 0.300 4.340 0.540 ;
        RECT  5.180 0.300 5.340 1.780 ;
        RECT  5.180 0.900 6.510 1.100 ;
        RECT  5.180 0.900 5.360 1.780 ;
        RECT  4.100 1.560 5.360 1.780 ;
        RECT  6.670 0.480 6.870 1.600 ;
        RECT  5.910 1.380 6.870 1.600 ;
        RECT  0.660 0.370 0.860 0.870 ;
        RECT  0.660 0.710 1.500 0.870 ;
        RECT  7.460 1.120 9.500 1.280 ;
        RECT  1.340 0.710 1.500 1.680 ;
        RECT  7.460 1.120 7.620 1.580 ;
        RECT  7.040 1.420 7.620 1.580 ;
        RECT  0.660 1.520 1.700 1.680 ;
        RECT  2.220 1.760 3.580 1.920 ;
        RECT  7.040 1.420 7.200 1.920 ;
        RECT  5.810 1.760 7.200 1.920 ;
        RECT  1.540 1.520 1.700 2.100 ;
        RECT  3.420 1.760 3.580 2.100 ;
        RECT  0.660 1.520 0.860 2.070 ;
        RECT  2.220 1.760 2.380 2.100 ;
        RECT  1.540 1.940 2.380 2.100 ;
        RECT  5.810 1.760 5.970 2.100 ;
        RECT  3.420 1.940 5.970 2.100 ;
        RECT  7.060 0.800 9.920 0.960 ;
        RECT  9.700 0.800 9.920 1.110 ;
        RECT  7.060 0.800 7.260 1.180 ;
        LAYER VTPH ;
        RECT  2.200 1.080 4.040 2.400 ;
        RECT  6.320 1.060 7.290 2.400 ;
        RECT  0.000 1.140 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.060 ;
        RECT  0.000 0.000 6.320 1.080 ;
        RECT  0.000 0.000 2.200 1.140 ;
        RECT  4.040 0.000 6.320 1.140 ;
        RECT  7.290 0.000 10.400 1.140 ;
    END
END LAGCEM6HM

MACRO LAGCEM4HM
    CLASS CORE ;
    FOREIGN LAGCEM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        ANTENNAGATEAREA 0.142  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.571  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.810 1.050 2.010 1.250 ;
        LAYER ME2 ;
        RECT  1.680 0.840 2.010 1.560 ;
        LAYER ME1 ;
        RECT  1.660 1.030 2.140 1.250 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.802  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.230 1.110 0.430 1.310 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.430 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.070 0.560 1.360 ;
        END
    END CK
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.412  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.940 1.580 7.100 1.740 ;
        RECT  6.900 0.480 7.100 1.740 ;
        RECT  5.580 0.480 7.100 0.640 ;
        RECT  5.940 1.580 6.140 2.100 ;
        RECT  5.580 0.320 5.780 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.740 1.900 7.020 2.540 ;
        RECT  5.080 1.800 5.240 2.540 ;
        RECT  3.960 2.080 4.240 2.540 ;
        RECT  1.980 1.800 2.140 2.540 ;
        RECT  0.640 1.840 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.140 -0.140 6.420 0.320 ;
        RECT  5.060 -0.140 5.260 0.600 ;
        RECT  3.560 -0.140 3.760 0.610 ;
        RECT  1.760 -0.140 2.040 0.540 ;
        RECT  0.660 -0.140 0.860 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.710 2.460 0.870 ;
        RECT  2.300 0.710 2.460 1.210 ;
        RECT  2.300 0.930 2.960 1.210 ;
        RECT  1.340 0.310 1.500 1.780 ;
        RECT  2.600 0.370 3.280 0.570 ;
        RECT  3.120 0.880 4.240 1.080 ;
        RECT  3.120 0.370 3.280 1.780 ;
        RECT  2.860 1.500 3.280 1.780 ;
        RECT  4.440 0.440 4.600 1.600 ;
        RECT  3.830 1.400 4.600 1.600 ;
        RECT  4.760 0.800 6.000 0.960 ;
        RECT  5.720 0.800 6.000 1.060 ;
        RECT  4.760 0.800 4.960 1.180 ;
        RECT  0.140 0.390 0.340 0.880 ;
        RECT  0.140 0.720 0.980 0.880 ;
        RECT  5.200 1.260 6.680 1.420 ;
        RECT  6.400 0.800 6.680 1.420 ;
        RECT  0.820 0.720 0.980 1.680 ;
        RECT  1.660 1.410 2.480 1.570 ;
        RECT  5.200 1.120 5.480 1.580 ;
        RECT  4.760 1.420 5.480 1.580 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  4.760 1.420 4.920 1.920 ;
        RECT  3.440 1.760 4.920 1.920 ;
        RECT  1.020 1.520 1.180 2.100 ;
        RECT  2.320 1.410 2.480 2.100 ;
        RECT  0.140 1.520 0.340 2.080 ;
        RECT  1.660 1.410 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  3.440 1.760 3.600 2.100 ;
        RECT  2.320 1.940 3.600 2.100 ;
        LAYER VTPH ;
        RECT  4.070 1.060 5.070 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.060 ;
        RECT  0.000 0.000 4.070 1.140 ;
        RECT  5.070 0.000 7.200 1.140 ;
    END
END LAGCEM4HM

MACRO LAGCEM3HM
    CLASS CORE ;
    FOREIGN LAGCEM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        ANTENNAGATEAREA 0.114  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.193  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.810 1.050 2.010 1.250 ;
        LAYER ME2 ;
        RECT  1.680 0.840 2.010 1.560 ;
        LAYER ME1 ;
        RECT  1.660 1.030 2.140 1.250 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        ANTENNAGATEAREA 0.118  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.316  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.230 1.110 0.430 1.310 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.430 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.070 0.560 1.360 ;
        END
    END CK
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.320  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.940 1.580 7.100 1.740 ;
        RECT  6.900 0.480 7.100 1.740 ;
        RECT  5.580 0.480 7.100 0.640 ;
        RECT  5.940 1.580 6.140 2.100 ;
        RECT  5.580 0.320 5.780 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.740 1.900 7.020 2.540 ;
        RECT  5.080 1.800 5.240 2.540 ;
        RECT  3.960 2.080 4.240 2.540 ;
        RECT  1.980 1.830 2.180 2.540 ;
        RECT  0.640 1.840 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.140 -0.140 6.420 0.320 ;
        RECT  5.060 -0.140 5.260 0.600 ;
        RECT  3.560 -0.140 3.760 0.610 ;
        RECT  1.760 -0.140 2.040 0.540 ;
        RECT  0.660 -0.140 0.860 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.340 0.710 2.960 0.870 ;
        RECT  2.760 0.710 2.960 1.210 ;
        RECT  1.340 0.310 1.500 1.780 ;
        RECT  2.550 0.380 3.280 0.540 ;
        RECT  3.120 0.880 4.240 1.080 ;
        RECT  3.120 0.380 3.280 1.780 ;
        RECT  2.860 1.500 3.280 1.780 ;
        RECT  4.440 0.440 4.600 1.600 ;
        RECT  3.830 1.400 4.600 1.600 ;
        RECT  4.760 0.800 6.000 0.960 ;
        RECT  5.720 0.800 6.000 1.060 ;
        RECT  4.760 0.800 4.960 1.180 ;
        RECT  0.140 0.390 0.340 0.880 ;
        RECT  0.140 0.720 0.980 0.880 ;
        RECT  5.200 1.260 6.680 1.420 ;
        RECT  6.400 0.800 6.680 1.420 ;
        RECT  0.820 0.720 0.980 1.680 ;
        RECT  1.660 1.410 2.560 1.570 ;
        RECT  5.200 1.120 5.480 1.580 ;
        RECT  4.760 1.420 5.480 1.580 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  4.760 1.420 4.920 1.920 ;
        RECT  3.440 1.760 4.920 1.920 ;
        RECT  1.020 1.520 1.180 2.100 ;
        RECT  2.400 1.410 2.560 2.100 ;
        RECT  0.140 1.520 0.340 2.080 ;
        RECT  1.660 1.410 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  3.440 1.760 3.600 2.100 ;
        RECT  2.400 1.940 3.600 2.100 ;
        LAYER VTPH ;
        RECT  4.070 1.060 5.070 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.060 ;
        RECT  0.000 0.000 4.070 1.140 ;
        RECT  5.070 0.000 7.200 1.140 ;
    END
END LAGCEM3HM

MACRO LAGCEM2HM
    CLASS CORE ;
    FOREIGN LAGCEM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        ANTENNAGATEAREA 0.092  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.446  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.040 0.300 1.240 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.980 0.560 1.310 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.297  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.720 1.040 1.920 1.240 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.920 1.560 ;
        LAYER ME1 ;
        RECT  1.660 1.040 2.310 1.320 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.352  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 1.440 6.600 2.080 ;
        RECT  6.400 0.480 6.600 2.080 ;
        RECT  5.860 0.480 6.600 0.640 ;
        RECT  5.860 0.320 6.060 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.280 1.750 5.480 2.540 ;
        RECT  4.000 2.080 4.280 2.540 ;
        RECT  1.980 1.800 2.140 2.540 ;
        RECT  0.660 1.830 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.420 -0.140 6.700 0.320 ;
        RECT  5.260 -0.140 5.460 0.600 ;
        RECT  4.040 -0.140 4.240 0.600 ;
        RECT  1.850 -0.140 2.130 0.540 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.220 0.300 1.500 0.560 ;
        RECT  1.340 0.720 2.840 0.880 ;
        RECT  2.680 0.720 2.840 1.310 ;
        RECT  1.340 0.300 1.500 1.780 ;
        RECT  2.800 0.360 3.160 0.560 ;
        RECT  3.000 0.900 4.380 1.100 ;
        RECT  3.000 0.360 3.160 1.780 ;
        RECT  2.760 1.620 3.160 1.780 ;
        RECT  3.740 1.400 4.780 1.560 ;
        RECT  4.540 0.320 4.780 1.600 ;
        RECT  4.500 1.400 4.780 1.600 ;
        RECT  0.100 0.350 0.380 0.820 ;
        RECT  0.100 0.660 0.980 0.820 ;
        RECT  0.820 0.660 0.980 1.640 ;
        RECT  5.400 1.120 5.680 1.560 ;
        RECT  4.940 1.400 5.680 1.560 ;
        RECT  0.140 1.480 1.180 1.640 ;
        RECT  1.660 1.480 2.480 1.640 ;
        RECT  4.940 1.400 5.100 1.920 ;
        RECT  3.350 1.760 5.100 1.920 ;
        RECT  1.020 1.480 1.180 2.100 ;
        RECT  2.320 1.480 2.480 2.100 ;
        RECT  0.140 1.480 0.340 2.030 ;
        RECT  1.660 1.480 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  3.350 1.420 3.510 2.100 ;
        RECT  2.320 1.940 3.510 2.100 ;
        RECT  4.960 0.800 6.240 0.960 ;
        RECT  4.960 0.800 5.160 1.140 ;
        LAYER VTPH ;
        RECT  4.000 1.070 4.980 2.400 ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.070 ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  4.980 0.000 6.800 1.140 ;
    END
END LAGCEM2HM

MACRO LAGCEM20HM
    CLASS CORE ;
    FOREIGN LAGCEM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.632  LAYER ME1  ;
        ANTENNAGATEAREA 0.632  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.891  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 0.980 2.300 1.180 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.560 ;
        LAYER ME1 ;
        RECT  0.440 0.980 2.520 1.200 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.708  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.040 0.480 4.540 0.860 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.520 1.500 21.500 1.660 ;
        RECT  21.340 0.480 21.500 1.660 ;
        RECT  13.000 0.480 21.500 0.640 ;
        RECT  20.280 1.500 20.560 2.100 ;
        RECT  18.960 0.320 19.160 0.640 ;
        RECT  18.600 1.500 18.880 2.100 ;
        RECT  17.280 0.330 17.480 0.640 ;
        RECT  16.840 1.500 17.200 2.100 ;
        RECT  15.420 0.330 15.620 0.640 ;
        RECT  15.240 1.500 15.520 2.100 ;
        RECT  14.120 0.330 14.320 0.640 ;
        RECT  13.520 1.500 13.800 2.100 ;
        RECT  13.000 0.330 13.200 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 21.600 2.540 ;
        RECT  21.120 1.880 21.400 2.540 ;
        RECT  19.440 1.900 19.720 2.540 ;
        RECT  17.760 1.900 18.040 2.540 ;
        RECT  16.080 1.900 16.360 2.540 ;
        RECT  14.400 1.900 14.680 2.540 ;
        RECT  12.680 1.820 12.880 2.540 ;
        RECT  11.020 2.080 11.300 2.540 ;
        RECT  6.520 2.080 6.800 2.540 ;
        RECT  5.320 2.080 5.600 2.540 ;
        RECT  4.120 2.080 4.400 2.540 ;
        RECT  2.740 1.830 2.940 2.540 ;
        RECT  1.700 1.830 1.900 2.540 ;
        RECT  0.660 1.830 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 21.600 0.140 ;
        RECT  19.480 -0.140 19.760 0.320 ;
        RECT  17.870 -0.140 18.570 0.320 ;
        RECT  16.170 -0.140 16.810 0.320 ;
        RECT  14.680 -0.140 14.960 0.320 ;
        RECT  13.520 -0.140 13.800 0.320 ;
        RECT  12.460 -0.140 12.760 0.630 ;
        RECT  10.900 -0.140 11.100 0.690 ;
        RECT  6.540 -0.140 6.820 0.510 ;
        RECT  5.500 -0.140 5.780 0.510 ;
        RECT  4.270 -0.140 4.550 0.320 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.680 1.440 7.450 1.600 ;
        RECT  5.020 0.410 5.220 0.860 ;
        RECT  6.060 0.410 6.260 0.860 ;
        RECT  7.120 0.410 7.320 0.860 ;
        RECT  8.240 0.620 8.520 0.860 ;
        RECT  9.320 0.620 9.600 0.860 ;
        RECT  5.020 0.700 9.600 0.860 ;
        RECT  3.420 1.020 10.220 1.180 ;
        RECT  9.900 0.960 10.220 1.240 ;
        RECT  3.420 0.320 3.700 1.600 ;
        RECT  11.670 0.620 11.980 1.390 ;
        RECT  11.140 1.190 11.980 1.390 ;
        RECT  11.780 0.620 11.980 1.780 ;
        RECT  7.680 0.300 9.960 0.460 ;
        RECT  11.270 0.300 12.300 0.460 ;
        RECT  9.800 0.300 9.960 0.680 ;
        RECT  7.680 0.300 7.960 0.540 ;
        RECT  8.800 0.300 9.080 0.540 ;
        RECT  9.800 0.520 10.540 0.680 ;
        RECT  12.140 0.300 12.300 1.280 ;
        RECT  12.140 0.800 20.780 0.960 ;
        RECT  11.270 0.300 11.430 1.030 ;
        RECT  10.380 0.870 11.430 1.030 ;
        RECT  12.140 0.800 12.360 1.280 ;
        RECT  10.380 0.520 10.540 1.560 ;
        RECT  9.920 1.400 10.540 1.560 ;
        RECT  9.920 1.400 10.200 1.780 ;
        RECT  7.640 1.620 10.200 1.780 ;
        RECT  0.140 0.340 0.340 0.820 ;
        RECT  1.180 0.340 1.380 0.820 ;
        RECT  2.220 0.340 2.420 0.820 ;
        RECT  0.140 0.660 3.060 0.820 ;
        RECT  20.980 1.000 21.180 1.280 ;
        RECT  12.560 1.120 21.180 1.280 ;
        RECT  2.900 0.660 3.060 1.670 ;
        RECT  12.560 1.120 12.720 1.640 ;
        RECT  12.360 1.480 12.720 1.640 ;
        RECT  0.140 1.510 3.260 1.670 ;
        RECT  3.100 1.510 3.260 1.920 ;
        RECT  3.100 1.760 7.120 1.920 ;
        RECT  10.480 1.760 11.620 1.920 ;
        RECT  6.960 1.760 7.120 2.100 ;
        RECT  11.460 1.760 11.620 2.100 ;
        RECT  0.140 1.510 0.340 1.970 ;
        RECT  1.180 1.510 1.380 1.990 ;
        RECT  2.220 1.510 2.420 1.990 ;
        RECT  10.480 1.760 10.640 2.100 ;
        RECT  6.960 1.940 10.640 2.100 ;
        RECT  12.360 1.480 12.520 2.100 ;
        RECT  11.460 1.940 12.520 2.100 ;
        LAYER VTPH ;
        RECT  3.240 1.080 7.630 2.400 ;
        RECT  0.000 1.140 21.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 21.600 1.080 ;
        RECT  0.000 0.000 3.240 1.140 ;
        RECT  7.630 0.000 21.600 1.140 ;
    END
END LAGCEM20HM

MACRO LAGCEM16HM
    CLASS CORE ;
    FOREIGN LAGCEM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.506  LAYER ME1  ;
        ANTENNAGATEAREA 0.506  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.992  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 0.980 1.500 1.180 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.280 0.980 2.000 1.200 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.566  LAYER ME2  ;
        ANTENNAGATEAREA 0.566  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 0.725  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.340 0.480 3.540 0.680 ;
        LAYER ME2 ;
        RECT  3.300 0.420 3.540 1.160 ;
        LAYER ME1 ;
        RECT  3.340 0.300 3.570 0.860 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.038  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.260 1.500 18.560 1.660 ;
        RECT  18.400 0.480 18.560 1.660 ;
        RECT  11.740 0.480 18.560 0.640 ;
        RECT  17.700 0.320 17.900 0.640 ;
        RECT  17.340 1.500 17.620 2.100 ;
        RECT  16.320 0.330 16.520 0.640 ;
        RECT  15.580 1.500 16.020 2.100 ;
        RECT  14.160 0.330 14.360 0.640 ;
        RECT  13.980 1.500 14.260 2.100 ;
        RECT  12.860 0.330 13.060 0.640 ;
        RECT  12.260 1.500 12.540 2.100 ;
        RECT  11.740 0.330 11.940 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.800 2.540 ;
        RECT  18.180 1.880 18.460 2.540 ;
        RECT  16.500 1.900 16.780 2.540 ;
        RECT  14.820 1.900 15.100 2.540 ;
        RECT  13.140 1.900 13.420 2.540 ;
        RECT  11.420 1.820 11.620 2.540 ;
        RECT  9.760 2.080 10.040 2.540 ;
        RECT  5.260 2.080 5.540 2.540 ;
        RECT  4.060 2.080 4.340 2.540 ;
        RECT  2.220 1.830 2.420 2.540 ;
        RECT  1.180 1.830 1.380 2.540 ;
        RECT  0.140 1.830 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.800 0.140 ;
        RECT  17.000 -0.140 17.310 0.320 ;
        RECT  14.910 -0.140 15.550 0.320 ;
        RECT  13.420 -0.140 13.700 0.320 ;
        RECT  12.260 -0.140 12.540 0.320 ;
        RECT  11.200 -0.140 11.500 0.630 ;
        RECT  9.640 -0.140 9.840 0.690 ;
        RECT  5.280 -0.140 5.560 0.510 ;
        RECT  4.240 -0.140 4.520 0.510 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.100 -0.140 0.380 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.420 1.440 6.190 1.600 ;
        RECT  3.760 0.410 3.960 0.860 ;
        RECT  4.800 0.410 5.000 0.860 ;
        RECT  5.860 0.410 6.060 0.860 ;
        RECT  6.980 0.620 7.260 0.860 ;
        RECT  8.060 0.620 8.340 0.860 ;
        RECT  3.760 0.700 8.340 0.860 ;
        RECT  2.900 1.020 8.960 1.180 ;
        RECT  8.640 0.960 8.960 1.240 ;
        RECT  2.900 0.320 3.180 1.680 ;
        RECT  10.410 0.620 10.720 1.390 ;
        RECT  9.880 1.190 10.720 1.390 ;
        RECT  10.520 0.620 10.720 1.780 ;
        RECT  6.420 0.300 8.700 0.460 ;
        RECT  10.010 0.300 11.040 0.460 ;
        RECT  8.540 0.300 8.700 0.680 ;
        RECT  6.420 0.300 6.700 0.540 ;
        RECT  7.540 0.300 7.820 0.540 ;
        RECT  8.540 0.520 9.280 0.680 ;
        RECT  10.880 0.300 11.040 1.280 ;
        RECT  10.880 0.800 17.850 0.960 ;
        RECT  10.010 0.300 10.170 1.030 ;
        RECT  9.120 0.870 10.170 1.030 ;
        RECT  10.880 0.800 11.100 1.280 ;
        RECT  9.120 0.520 9.280 1.560 ;
        RECT  8.660 1.400 9.280 1.560 ;
        RECT  8.660 1.400 8.940 1.780 ;
        RECT  6.380 1.620 8.940 1.780 ;
        RECT  0.660 0.340 0.860 0.820 ;
        RECT  1.700 0.340 1.900 0.820 ;
        RECT  0.660 0.660 2.540 0.820 ;
        RECT  18.040 1.000 18.240 1.280 ;
        RECT  11.300 1.120 18.240 1.280 ;
        RECT  2.380 0.660 2.540 1.670 ;
        RECT  11.300 1.120 11.460 1.640 ;
        RECT  11.100 1.480 11.460 1.640 ;
        RECT  0.660 1.510 2.740 1.670 ;
        RECT  3.600 1.760 5.860 1.920 ;
        RECT  9.220 1.760 10.360 1.920 ;
        RECT  2.580 1.510 2.740 2.100 ;
        RECT  5.700 1.760 5.860 2.100 ;
        RECT  10.200 1.760 10.360 2.100 ;
        RECT  0.660 1.510 0.860 1.990 ;
        RECT  1.700 1.510 1.900 1.990 ;
        RECT  3.600 1.760 3.760 2.100 ;
        RECT  2.580 1.940 3.760 2.100 ;
        RECT  9.220 1.760 9.380 2.100 ;
        RECT  5.700 1.940 9.380 2.100 ;
        RECT  11.100 1.480 11.260 2.100 ;
        RECT  10.200 1.940 11.260 2.100 ;
        LAYER VTPH ;
        RECT  3.240 1.080 6.370 2.400 ;
        RECT  0.000 1.140 18.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.800 1.080 ;
        RECT  0.000 0.000 3.240 1.140 ;
        RECT  6.370 0.000 18.800 1.140 ;
    END
END LAGCEM16HM

MACRO LAGCEM12HM
    CLASS CORE ;
    FOREIGN LAGCEM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.388  LAYER ME1  ;
        ANTENNAGATEAREA 0.388  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.690  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 0.980 1.100 1.180 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.440 0.980 1.480 1.200 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.425  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 0.300 3.140 0.860 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.499  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.280 1.500 15.900 1.660 ;
        RECT  15.740 0.480 15.900 1.660 ;
        RECT  10.760 0.480 15.900 0.640 ;
        RECT  15.040 0.350 15.320 0.640 ;
        RECT  14.680 1.500 15.100 2.100 ;
        RECT  13.180 0.330 13.380 0.640 ;
        RECT  13.000 1.500 13.280 2.100 ;
        RECT  11.880 0.330 12.080 0.640 ;
        RECT  11.280 1.500 11.560 2.100 ;
        RECT  10.760 0.330 10.960 0.640 ;
        END
    END GCK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.000 2.540 ;
        RECT  15.520 1.880 15.800 2.540 ;
        RECT  13.840 1.900 14.120 2.540 ;
        RECT  12.160 1.900 12.440 2.540 ;
        RECT  10.440 1.820 10.640 2.540 ;
        RECT  8.780 2.080 9.060 2.540 ;
        RECT  4.280 2.080 4.560 2.540 ;
        RECT  3.080 2.080 3.360 2.540 ;
        RECT  1.700 1.830 1.900 2.540 ;
        RECT  0.660 1.830 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.000 0.140 ;
        RECT  13.930 -0.140 14.570 0.320 ;
        RECT  12.440 -0.140 12.720 0.320 ;
        RECT  11.280 -0.140 11.560 0.320 ;
        RECT  10.220 -0.140 10.520 0.630 ;
        RECT  8.660 -0.140 8.860 0.690 ;
        RECT  4.300 -0.140 4.580 0.510 ;
        RECT  3.300 -0.140 3.540 0.630 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.560 1.440 5.210 1.600 ;
        RECT  3.820 0.410 4.020 0.860 ;
        RECT  4.880 0.410 5.080 0.860 ;
        RECT  6.000 0.620 6.280 0.860 ;
        RECT  7.080 0.620 7.360 0.860 ;
        RECT  3.820 0.700 7.360 0.860 ;
        RECT  2.380 0.320 2.660 1.180 ;
        RECT  2.380 1.020 7.980 1.180 ;
        RECT  7.660 0.960 7.980 1.240 ;
        RECT  2.380 0.320 2.580 1.740 ;
        RECT  9.430 0.620 9.740 1.390 ;
        RECT  8.900 1.190 9.740 1.390 ;
        RECT  9.540 0.620 9.740 1.780 ;
        RECT  5.440 0.300 7.720 0.460 ;
        RECT  9.030 0.300 10.060 0.460 ;
        RECT  7.560 0.300 7.720 0.680 ;
        RECT  5.440 0.300 5.720 0.540 ;
        RECT  6.560 0.300 6.840 0.540 ;
        RECT  7.560 0.520 8.300 0.680 ;
        RECT  9.900 0.300 10.060 1.280 ;
        RECT  9.900 0.800 15.180 0.960 ;
        RECT  9.030 0.300 9.190 1.030 ;
        RECT  8.140 0.870 9.190 1.030 ;
        RECT  9.900 0.800 10.120 1.280 ;
        RECT  8.140 0.520 8.300 1.560 ;
        RECT  7.680 1.400 8.300 1.560 ;
        RECT  7.680 1.400 7.960 1.780 ;
        RECT  5.400 1.620 7.960 1.780 ;
        RECT  0.140 0.340 0.340 0.820 ;
        RECT  1.180 0.340 1.380 0.820 ;
        RECT  0.140 0.660 2.020 0.820 ;
        RECT  15.380 1.000 15.580 1.280 ;
        RECT  10.320 1.120 15.580 1.280 ;
        RECT  1.860 0.660 2.020 1.670 ;
        RECT  10.320 1.120 10.480 1.640 ;
        RECT  10.120 1.480 10.480 1.640 ;
        RECT  0.140 1.510 2.220 1.670 ;
        RECT  2.760 1.760 4.880 1.920 ;
        RECT  8.240 1.760 9.380 1.920 ;
        RECT  2.060 1.510 2.220 2.100 ;
        RECT  4.720 1.760 4.880 2.100 ;
        RECT  9.220 1.760 9.380 2.100 ;
        RECT  0.140 1.510 0.340 1.990 ;
        RECT  1.180 1.510 1.380 1.990 ;
        RECT  2.760 1.760 2.920 2.100 ;
        RECT  2.060 1.940 2.920 2.100 ;
        RECT  8.240 1.760 8.400 2.100 ;
        RECT  4.720 1.940 8.400 2.100 ;
        RECT  10.120 1.480 10.280 2.100 ;
        RECT  9.220 1.940 10.280 2.100 ;
        LAYER VTPH ;
        RECT  2.800 1.080 5.390 2.400 ;
        RECT  0.000 1.140 16.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.000 1.080 ;
        RECT  0.000 0.000 2.800 1.140 ;
        RECT  5.390 0.000 16.000 1.140 ;
    END
END LAGCEM12HM

MACRO LAGCECSM8HM
    CLASS CORE ;
    FOREIGN LAGCECSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.361  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.000 1.245 8.750 1.405 ;
        RECT  8.395 1.120 8.750 1.405 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.245 7.160 2.100 ;
        RECT  6.255 1.300 6.415 2.100 ;
        RECT  5.560 1.300 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.817  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.165 0.430 11.495 0.710 ;
        RECT  11.120 0.660 11.340 2.100 ;
        RECT  10.080 1.410 11.340 1.675 ;
        RECT  10.160 0.660 11.340 0.820 ;
        RECT  10.160 0.325 10.380 0.820 ;
        RECT  10.080 1.410 10.300 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  11.580 1.440 11.860 2.540 ;
        RECT  10.540 1.835 10.820 2.540 ;
        RECT  9.500 1.900 9.780 2.540 ;
        RECT  7.340 1.765 7.620 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  10.620 -0.140 10.900 0.500 ;
        RECT  9.540 -0.140 9.820 0.320 ;
        RECT  8.420 -0.140 8.700 0.320 ;
        RECT  7.340 -0.140 7.620 0.500 ;
        RECT  6.320 -0.140 6.480 0.935 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.785 0.800 6.060 1.140 ;
        RECT  5.220 0.955 6.060 1.140 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.680 0.660 7.680 0.850 ;
        RECT  7.520 0.800 9.440 0.960 ;
        RECT  7.520 0.800 7.800 1.050 ;
        RECT  9.160 0.800 9.440 1.140 ;
        RECT  6.680 0.660 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.840 0.400 8.170 0.640 ;
        RECT  8.970 0.370 9.265 0.640 ;
        RECT  7.840 0.480 9.900 0.640 ;
        RECT  9.740 1.020 10.715 1.180 ;
        RECT  9.180 1.580 9.900 1.740 ;
        RECT  9.740 0.480 9.900 1.740 ;
        RECT  8.395 1.735 9.340 1.895 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.220 12.000 2.400 ;
        RECT  7.260 1.140 12.000 2.400 ;
        RECT  0.000 1.320 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.140 ;
        RECT  4.220 0.000 7.260 1.220 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM8HM

MACRO LAGCECSM6HM
    CLASS CORE ;
    FOREIGN LAGCECSM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.294  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.000 1.190 8.720 1.560 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.190 7.160 2.100 ;
        RECT  6.255 1.350 6.415 2.100 ;
        RECT  5.560 1.350 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.692  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.120 1.015 11.340 2.100 ;
        RECT  10.080 1.015 11.340 1.235 ;
        RECT  10.080 0.325 10.325 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.540 1.440 10.820 2.540 ;
        RECT  9.500 1.900 9.780 2.540 ;
        RECT  7.340 1.900 7.620 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.660 -0.140 10.940 0.620 ;
        RECT  9.540 -0.140 9.820 0.320 ;
        RECT  8.420 -0.140 8.700 0.320 ;
        RECT  7.340 -0.140 7.620 0.620 ;
        RECT  6.320 -0.140 6.480 0.935 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.220 0.955 6.060 1.190 ;
        RECT  5.785 0.800 6.060 1.190 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.680 0.590 7.060 1.030 ;
        RECT  6.680 0.820 9.570 1.030 ;
        RECT  6.680 0.590 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.840 0.400 8.170 0.660 ;
        RECT  8.970 0.385 9.275 0.660 ;
        RECT  7.840 0.500 9.900 0.660 ;
        RECT  9.160 1.580 9.900 1.740 ;
        RECT  9.740 0.500 9.900 1.740 ;
        RECT  8.480 1.735 9.320 1.895 ;
        RECT  8.480 1.735 8.640 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.210 11.600 2.400 ;
        RECT  8.640 1.140 11.600 2.400 ;
        RECT  0.000 1.320 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.140 ;
        RECT  4.220 0.000 8.640 1.210 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM6HM

MACRO LAGCECSM4HM
    CLASS CORE ;
    FOREIGN LAGCECSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.215  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.000 1.190 7.880 1.420 ;
        RECT  7.000 1.190 7.560 1.560 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.190 7.160 2.100 ;
        RECT  6.255 1.350 6.415 2.100 ;
        RECT  5.560 1.350 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.880 0.325 9.120 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.340 1.440 9.620 2.540 ;
        RECT  8.300 1.900 8.580 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.420 -0.140 9.700 0.650 ;
        RECT  8.340 -0.140 8.620 0.320 ;
        RECT  7.320 -0.140 7.540 0.650 ;
        RECT  6.320 -0.140 6.480 0.935 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.220 0.955 6.060 1.190 ;
        RECT  5.785 0.800 6.060 1.190 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.680 0.590 7.060 1.030 ;
        RECT  6.680 0.820 8.280 1.030 ;
        RECT  6.680 0.590 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.840 0.300 8.000 0.645 ;
        RECT  7.840 0.485 8.700 0.645 ;
        RECT  7.960 1.580 8.700 1.740 ;
        RECT  8.540 0.485 8.700 1.740 ;
        RECT  7.320 1.735 8.120 1.895 ;
        RECT  7.320 1.735 7.480 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.210 10.000 2.400 ;
        RECT  7.480 1.140 10.000 2.400 ;
        RECT  0.000 1.320 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  4.220 0.000 7.480 1.210 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM4HM

MACRO LAGCECSM3HM
    CLASS CORE ;
    FOREIGN LAGCECSM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.215  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.000 1.190 7.785 1.420 ;
        RECT  7.000 1.190 7.560 1.560 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.190 7.160 2.100 ;
        RECT  6.255 1.350 6.415 2.100 ;
        RECT  5.560 1.350 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.354  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.880 0.325 9.120 2.040 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.340 1.600 9.620 2.540 ;
        RECT  8.300 1.900 8.580 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  8.340 -0.140 8.620 0.360 ;
        RECT  7.020 -0.140 7.315 0.550 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.220 0.955 6.060 1.190 ;
        RECT  5.785 0.800 6.060 1.190 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.320 0.640 6.840 0.920 ;
        RECT  6.680 0.840 8.280 1.000 ;
        RECT  7.945 0.840 8.280 1.040 ;
        RECT  6.680 0.640 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.840 0.300 8.000 0.680 ;
        RECT  7.840 0.520 8.700 0.680 ;
        RECT  7.960 1.580 8.700 1.740 ;
        RECT  8.540 0.520 8.700 1.740 ;
        RECT  7.320 1.735 8.120 1.895 ;
        RECT  7.320 1.735 7.480 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.210 10.000 2.400 ;
        RECT  7.480 1.140 10.000 2.400 ;
        RECT  0.000 1.320 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  4.220 0.000 7.480 1.210 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM3HM

MACRO LAGCECSM2HM
    CLASS CORE ;
    FOREIGN LAGCECSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.205  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.000 1.220 7.810 1.420 ;
        RECT  7.000 1.220 7.560 1.560 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.220 7.160 2.100 ;
        RECT  6.255 1.350 6.415 2.100 ;
        RECT  5.560 1.350 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.326  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.880 0.325 9.100 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.300 1.900 8.580 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.250 -0.140 8.530 0.320 ;
        RECT  7.020 -0.140 7.315 0.550 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.540 1.180 3.870 1.340 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.220 0.955 6.010 1.190 ;
        RECT  5.735 0.800 6.010 1.190 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.970 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.150 0.640 ;
        RECT  4.860 0.480 6.150 0.640 ;
        RECT  3.970 0.380 4.200 1.020 ;
        RECT  2.975 0.840 4.200 1.020 ;
        RECT  2.975 0.840 3.255 1.060 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.320 0.640 6.735 0.920 ;
        RECT  6.575 0.820 8.320 1.040 ;
        RECT  6.575 0.640 6.735 1.780 ;
        RECT  6.575 1.520 6.840 1.780 ;
        RECT  7.680 0.300 7.840 0.640 ;
        RECT  7.680 0.480 8.700 0.640 ;
        RECT  7.960 1.580 8.700 1.740 ;
        RECT  8.540 0.480 8.700 1.740 ;
        RECT  7.320 1.735 8.120 1.895 ;
        RECT  7.320 1.735 7.480 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  6.295 1.220 9.200 2.400 ;
        RECT  7.480 1.140 9.200 2.400 ;
        RECT  0.000 1.320 9.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.200 1.140 ;
        RECT  4.220 0.000 7.480 1.220 ;
        RECT  4.220 0.000 6.295 1.320 ;
    END
END LAGCECSM2HM

MACRO LAGCECSM20HM
    CLASS CORE ;
    FOREIGN LAGCECSM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.768  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.295 1.435 11.955 1.595 ;
        RECT  11.675 1.120 11.955 1.595 ;
        RECT  7.000 1.330 10.575 1.500 ;
        RECT  9.530 1.120 9.810 1.500 ;
        RECT  7.600 1.120 7.950 1.500 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.330 7.160 2.100 ;
        RECT  6.255 1.300 6.415 2.100 ;
        RECT  5.560 1.300 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.942  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.420 0.900 17.640 2.100 ;
        RECT  15.400 0.900 17.640 1.265 ;
        RECT  16.380 0.900 16.600 2.100 ;
        RECT  15.560 0.335 15.860 1.265 ;
        RECT  15.400 0.665 15.620 2.100 ;
        RECT  13.320 1.340 15.620 1.660 ;
        RECT  13.560 0.665 15.860 0.860 ;
        RECT  14.520 0.335 14.820 0.860 ;
        RECT  14.360 1.340 14.580 2.100 ;
        RECT  13.560 0.325 13.780 0.860 ;
        RECT  13.320 1.340 13.540 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.400 2.540 ;
        RECT  17.940 1.440 18.220 2.540 ;
        RECT  16.900 1.440 17.180 2.540 ;
        RECT  15.860 1.440 16.140 2.540 ;
        RECT  14.820 1.820 15.100 2.540 ;
        RECT  13.780 1.820 14.060 2.540 ;
        RECT  12.740 1.900 13.020 2.540 ;
        RECT  10.620 2.080 10.900 2.540 ;
        RECT  8.460 2.080 8.740 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.400 0.140 ;
        RECT  16.100 -0.140 16.380 0.680 ;
        RECT  15.060 -0.140 15.340 0.505 ;
        RECT  14.020 -0.140 14.300 0.505 ;
        RECT  12.940 -0.140 13.220 0.320 ;
        RECT  11.820 -0.140 12.100 0.320 ;
        RECT  10.700 -0.140 10.980 0.320 ;
        RECT  9.580 -0.140 9.860 0.320 ;
        RECT  8.460 -0.140 8.740 0.320 ;
        RECT  7.335 -0.140 7.615 0.625 ;
        RECT  6.320 -0.140 6.480 0.875 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.785 0.800 6.060 1.140 ;
        RECT  5.220 0.955 6.060 1.140 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.680 0.530 7.060 0.960 ;
        RECT  6.680 0.800 12.840 0.960 ;
        RECT  10.675 0.800 10.955 1.110 ;
        RECT  12.560 0.800 12.840 1.110 ;
        RECT  8.430 0.800 8.755 1.140 ;
        RECT  6.680 0.530 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.865 0.400 8.195 0.640 ;
        RECT  8.985 0.400 9.315 0.640 ;
        RECT  10.105 0.400 10.435 0.640 ;
        RECT  7.865 0.480 13.160 0.640 ;
        RECT  13.000 1.020 14.960 1.180 ;
        RECT  13.000 0.480 13.160 1.740 ;
        RECT  12.415 1.580 13.160 1.740 ;
        RECT  12.415 1.580 12.575 1.915 ;
        RECT  7.345 1.755 12.575 1.915 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.220 18.400 2.400 ;
        RECT  7.070 1.140 18.400 2.400 ;
        RECT  0.000 1.320 18.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.400 1.140 ;
        RECT  4.220 0.000 7.070 1.220 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM20HM

MACRO LAGCECSM16HM
    CLASS CORE ;
    FOREIGN LAGCECSM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.632  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.000 1.330 10.920 1.500 ;
        RECT  10.620 1.120 10.920 1.500 ;
        RECT  8.470 1.120 8.750 1.500 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.330 7.160 2.100 ;
        RECT  6.255 1.300 6.415 2.100 ;
        RECT  5.560 1.300 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.320 0.930 15.540 2.100 ;
        RECT  14.340 0.930 15.540 1.265 ;
        RECT  14.420 0.335 14.720 0.665 ;
        RECT  14.340 0.665 14.640 1.265 ;
        RECT  14.340 0.665 14.560 2.100 ;
        RECT  12.260 1.340 14.560 1.660 ;
        RECT  12.420 0.665 14.640 0.860 ;
        RECT  13.380 0.335 13.680 0.860 ;
        RECT  13.300 1.340 13.520 2.100 ;
        RECT  12.420 0.325 12.640 0.860 ;
        RECT  12.260 1.340 12.480 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.400 2.540 ;
        RECT  15.840 1.440 16.120 2.540 ;
        RECT  14.800 1.440 15.080 2.540 ;
        RECT  13.760 1.820 14.040 2.540 ;
        RECT  12.720 1.820 13.000 2.540 ;
        RECT  11.680 1.900 11.960 2.540 ;
        RECT  9.560 2.080 9.840 2.540 ;
        RECT  7.400 1.755 7.680 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.400 0.140 ;
        RECT  13.920 -0.140 14.200 0.505 ;
        RECT  12.880 -0.140 13.160 0.505 ;
        RECT  11.800 -0.140 12.080 0.320 ;
        RECT  10.680 -0.140 10.960 0.320 ;
        RECT  9.560 -0.140 9.840 0.320 ;
        RECT  8.440 -0.140 8.720 0.320 ;
        RECT  7.320 -0.140 7.600 0.505 ;
        RECT  6.320 -0.140 6.480 0.875 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.785 0.800 6.060 1.140 ;
        RECT  5.220 0.955 6.060 1.140 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.680 0.530 7.060 0.960 ;
        RECT  6.680 0.800 11.700 0.960 ;
        RECT  9.545 0.800 9.865 1.050 ;
        RECT  7.615 0.800 7.900 1.110 ;
        RECT  11.420 0.800 11.700 1.135 ;
        RECT  6.680 0.530 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.845 0.400 8.175 0.640 ;
        RECT  8.965 0.400 9.295 0.640 ;
        RECT  7.845 0.480 12.080 0.640 ;
        RECT  11.920 1.020 13.900 1.180 ;
        RECT  11.920 0.480 12.080 1.740 ;
        RECT  11.355 1.580 12.080 1.740 ;
        RECT  11.355 1.580 11.515 1.915 ;
        RECT  8.450 1.755 11.515 1.915 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.220 16.400 2.400 ;
        RECT  7.070 1.140 16.400 2.400 ;
        RECT  0.000 1.320 16.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.400 1.140 ;
        RECT  4.220 0.000 7.070 1.220 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM16HM

MACRO LAGCECSM12HM
    CLASS CORE ;
    FOREIGN LAGCECSM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.497  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.810 1.435 9.735 1.595 ;
        RECT  9.390 1.120 9.735 1.595 ;
        RECT  7.000 1.330 8.010 1.500 ;
        RECT  7.460 1.120 7.740 1.500 ;
        RECT  6.255 1.940 7.160 2.100 ;
        RECT  7.000 1.330 7.160 2.100 ;
        RECT  6.255 1.300 6.415 2.100 ;
        RECT  5.560 1.300 6.415 1.510 ;
        END
    END CKB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.050 1.100 1.960 ;
        END
    END E
    PIN GCK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.140 0.900 13.360 2.100 ;
        RECT  12.100 0.900 13.360 1.265 ;
        RECT  12.180 0.335 12.480 1.265 ;
        RECT  12.100 0.665 12.320 2.100 ;
        RECT  11.060 1.340 12.320 1.660 ;
        RECT  11.220 0.665 12.480 0.860 ;
        RECT  11.220 0.325 11.440 0.860 ;
        RECT  11.060 1.340 11.280 2.100 ;
        END
    END GCK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.050 0.700 1.560 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.600 1.440 13.880 2.540 ;
        RECT  12.560 1.440 12.840 2.540 ;
        RECT  11.520 1.820 11.800 2.540 ;
        RECT  10.480 1.900 10.760 2.540 ;
        RECT  8.360 2.080 8.640 2.540 ;
        RECT  5.880 1.770 6.095 2.540 ;
        RECT  4.880 1.710 5.040 2.540 ;
        RECT  2.960 1.860 3.240 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  12.720 -0.140 13.000 0.650 ;
        RECT  11.680 -0.140 11.960 0.505 ;
        RECT  10.600 -0.140 10.880 0.320 ;
        RECT  9.480 -0.140 9.760 0.320 ;
        RECT  8.360 -0.140 8.640 0.320 ;
        RECT  7.280 -0.140 7.560 0.500 ;
        RECT  6.320 -0.140 6.480 0.875 ;
        RECT  5.170 -0.140 5.450 0.320 ;
        RECT  3.135 -0.140 3.500 0.570 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.380 0.320 0.840 ;
        RECT  1.200 0.320 1.360 0.840 ;
        RECT  0.160 0.680 1.360 0.840 ;
        RECT  1.535 0.300 2.700 0.460 ;
        RECT  2.540 0.300 2.700 1.035 ;
        RECT  1.535 0.300 1.695 1.160 ;
        RECT  1.380 1.000 1.540 1.335 ;
        RECT  2.000 0.620 2.280 1.380 ;
        RECT  3.475 1.070 3.870 1.230 ;
        RECT  1.875 1.220 3.650 1.380 ;
        RECT  1.875 1.220 2.035 1.990 ;
        RECT  1.645 1.635 2.035 1.990 ;
        RECT  4.360 0.700 4.705 0.900 ;
        RECT  2.200 1.540 3.560 1.700 ;
        RECT  3.400 1.540 3.560 2.100 ;
        RECT  2.200 1.540 2.485 1.980 ;
        RECT  4.360 0.700 4.520 2.100 ;
        RECT  3.400 1.940 4.520 2.100 ;
        RECT  5.785 0.800 6.060 1.140 ;
        RECT  5.220 0.955 6.060 1.140 ;
        RECT  4.700 1.165 5.380 1.460 ;
        RECT  5.220 0.955 5.380 1.970 ;
        RECT  5.220 1.810 5.660 1.970 ;
        RECT  3.915 0.380 5.020 0.540 ;
        RECT  5.840 0.300 6.160 0.640 ;
        RECT  4.860 0.480 6.160 0.640 ;
        RECT  3.915 0.380 4.200 0.910 ;
        RECT  2.975 0.730 4.200 0.910 ;
        RECT  2.975 0.730 3.255 0.960 ;
        RECT  4.030 0.380 4.200 1.680 ;
        RECT  3.760 1.500 4.200 1.680 ;
        RECT  3.760 1.500 3.960 1.780 ;
        RECT  6.680 0.530 7.060 0.960 ;
        RECT  6.680 0.800 10.500 0.960 ;
        RECT  10.220 0.800 10.500 1.140 ;
        RECT  8.310 0.800 8.620 1.170 ;
        RECT  6.680 0.530 6.840 1.780 ;
        RECT  6.575 1.490 6.840 1.780 ;
        RECT  7.765 0.400 8.095 0.640 ;
        RECT  7.765 0.480 10.880 0.640 ;
        RECT  10.720 1.020 11.875 1.180 ;
        RECT  10.720 0.480 10.880 1.740 ;
        RECT  10.155 1.580 10.880 1.740 ;
        RECT  10.155 1.580 10.315 1.915 ;
        RECT  7.340 1.755 10.315 1.915 ;
        RECT  7.340 1.660 7.550 2.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.220 2.400 ;
        RECT  0.000 1.260 4.700 2.400 ;
        RECT  6.295 1.220 14.000 2.400 ;
        RECT  7.070 1.140 14.000 2.400 ;
        RECT  0.000 1.320 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.140 ;
        RECT  4.220 0.000 7.070 1.220 ;
        RECT  4.220 0.000 6.295 1.260 ;
        RECT  4.700 0.000 6.295 1.320 ;
    END
END LAGCECSM12HM

MACRO LACRSM4HM
    CLASS CORE ;
    FOREIGN LACRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        ANTENNAGATEAREA 0.092  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 22.342  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.620 0.700 4.330 0.920 ;
        RECT  4.110 0.620 4.330 0.920 ;
        RECT  2.620 0.300 2.780 0.920 ;
        RECT  1.060 0.300 2.780 0.500 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        ANTENNAGATEAREA 0.143  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.714  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.510 1.290 5.710 1.490 ;
        LAYER ME2 ;
        RECT  5.510 1.100 5.900 1.680 ;
        LAYER ME1 ;
        RECT  5.450 0.960 5.750 1.680 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.090  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 0.760 1.500 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.440 1.500 1.160 ;
        LAYER ME1 ;
        RECT  1.240 0.660 1.980 0.960 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.204  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 3.010 1.600 ;
        RECT  0.500 1.020 0.710 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.300 0.840 8.770 1.160 ;
        RECT  8.300 0.390 8.580 2.060 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.535  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.840 1.230 7.500 1.600 ;
        RECT  7.300 0.400 7.500 1.600 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  8.820 1.490 9.100 2.540 ;
        RECT  7.590 2.080 7.950 2.540 ;
        RECT  6.390 2.080 6.750 2.540 ;
        RECT  5.350 1.900 5.630 2.540 ;
        RECT  4.310 1.900 4.590 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.820 -0.140 9.100 0.670 ;
        RECT  7.780 -0.140 8.060 0.660 ;
        RECT  6.740 -0.140 7.020 0.680 ;
        RECT  4.810 -0.140 4.970 0.660 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.030 0.840 ;
        RECT  0.870 0.680 1.030 1.280 ;
        RECT  2.260 0.660 2.460 1.280 ;
        RECT  0.870 1.120 3.460 1.280 ;
        RECT  0.140 0.410 0.340 2.080 ;
        RECT  2.940 0.300 4.650 0.460 ;
        RECT  2.940 0.300 3.220 0.540 ;
        RECT  4.490 0.300 4.650 1.240 ;
        RECT  4.490 0.960 4.870 1.240 ;
        RECT  3.670 1.080 4.870 1.240 ;
        RECT  3.670 1.080 3.830 1.600 ;
        RECT  3.280 1.440 3.830 1.600 ;
        RECT  1.220 1.760 3.450 1.920 ;
        RECT  3.280 1.440 3.450 2.020 ;
        RECT  2.970 1.760 3.450 2.020 ;
        RECT  5.130 0.430 6.120 0.630 ;
        RECT  5.960 0.430 6.120 1.300 ;
        RECT  5.130 0.430 5.290 1.700 ;
        RECT  3.990 1.540 5.290 1.700 ;
        RECT  3.990 1.540 4.150 2.100 ;
        RECT  3.750 1.940 4.150 2.100 ;
        RECT  4.790 1.540 5.150 2.100 ;
        RECT  6.280 0.410 6.440 1.920 ;
        RECT  5.910 1.640 6.440 1.920 ;
        RECT  7.980 0.920 8.140 1.920 ;
        RECT  5.910 1.760 8.140 1.920 ;
        LAYER VTPH ;
        RECT  6.790 1.080 7.520 2.400 ;
        RECT  0.000 1.140 9.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.200 1.080 ;
        RECT  0.000 0.000 6.790 1.140 ;
        RECT  7.520 0.000 9.200 1.140 ;
    END
END LACRSM4HM

MACRO LACRSM2HM
    CLASS CORE ;
    FOREIGN LACRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.090  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 0.760 1.500 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.440 1.500 1.160 ;
        LAYER ME1 ;
        RECT  1.240 0.660 1.980 0.960 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        ANTENNAGATEAREA 0.143  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.714  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.510 1.290 5.710 1.490 ;
        LAYER ME2 ;
        RECT  5.300 1.230 5.900 1.570 ;
        LAYER ME1 ;
        RECT  5.450 0.960 5.750 1.680 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        ANTENNAGATEAREA 0.092  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 22.342  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.620 0.700 4.330 0.920 ;
        RECT  4.070 0.620 4.330 0.920 ;
        RECT  2.620 0.300 2.780 0.920 ;
        RECT  1.060 0.300 2.780 0.500 ;
        END
    END RB
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 3.010 1.600 ;
        RECT  0.500 1.020 0.710 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.300 0.390 8.700 2.060 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.840 1.240 7.500 1.600 ;
        RECT  7.300 0.400 7.500 1.600 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.740 2.080 8.020 2.540 ;
        RECT  6.430 2.080 6.710 2.540 ;
        RECT  5.350 1.900 5.630 2.540 ;
        RECT  4.310 1.900 4.590 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.780 -0.140 8.060 0.660 ;
        RECT  6.740 -0.140 7.020 0.720 ;
        RECT  4.810 -0.140 4.970 0.660 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.030 0.840 ;
        RECT  0.870 0.680 1.030 1.280 ;
        RECT  2.260 0.660 2.460 1.280 ;
        RECT  0.870 1.120 3.460 1.280 ;
        RECT  0.140 0.300 0.340 1.950 ;
        RECT  2.940 0.300 4.650 0.460 ;
        RECT  2.940 0.300 3.260 0.540 ;
        RECT  4.490 0.300 4.650 1.240 ;
        RECT  4.490 0.960 4.870 1.240 ;
        RECT  3.670 1.080 4.870 1.240 ;
        RECT  3.670 1.080 3.830 1.600 ;
        RECT  3.280 1.440 3.830 1.600 ;
        RECT  1.220 1.760 3.450 1.920 ;
        RECT  3.280 1.440 3.450 2.020 ;
        RECT  2.970 1.760 3.450 2.020 ;
        RECT  5.130 0.430 6.120 0.630 ;
        RECT  5.960 0.430 6.120 1.300 ;
        RECT  5.130 0.430 5.290 1.700 ;
        RECT  3.990 1.540 5.290 1.700 ;
        RECT  3.990 1.540 4.150 2.100 ;
        RECT  3.750 1.940 4.150 2.100 ;
        RECT  4.830 1.540 5.110 2.100 ;
        RECT  6.280 0.410 6.440 1.920 ;
        RECT  5.910 1.640 6.440 1.920 ;
        RECT  7.980 0.920 8.140 1.920 ;
        RECT  5.910 1.760 8.140 1.920 ;
        LAYER VTPH ;
        RECT  6.790 1.080 7.520 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.080 ;
        RECT  0.000 0.000 6.790 1.140 ;
        RECT  7.520 0.000 8.800 1.140 ;
    END
END LACRSM2HM

MACRO LACRSM1HM
    CLASS CORE ;
    FOREIGN LACRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.388  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.760 1.900 0.960 ;
        LAYER ME2 ;
        RECT  1.700 0.440 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.320 0.660 2.060 0.960 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        ANTENNAGATEAREA 0.104  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 15.241  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.590 1.260 0.790 1.460 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.790 1.680 ;
        LAYER ME1 ;
        RECT  0.580 1.440 3.060 1.600 ;
        RECT  0.580 1.020 0.790 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.340 0.390 8.700 1.790 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.332  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.070 1.240 7.580 1.600 ;
        RECT  7.380 0.400 7.580 1.600 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 26.880  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.700 0.700 4.410 0.920 ;
        RECT  4.150 0.620 4.410 0.920 ;
        RECT  2.700 0.300 2.860 0.920 ;
        RECT  1.140 0.300 2.860 0.500 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.262  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.580 1.290 5.780 1.490 ;
        LAYER ME2 ;
        RECT  5.300 1.230 5.900 1.570 ;
        LAYER ME1 ;
        RECT  5.530 0.960 5.830 1.680 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.780 2.080 8.060 2.540 ;
        RECT  6.510 2.080 6.790 2.540 ;
        RECT  5.430 1.880 5.710 2.540 ;
        RECT  4.390 1.880 4.670 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        RECT  0.740 2.080 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.820 -0.140 8.100 0.660 ;
        RECT  6.820 -0.140 7.100 0.720 ;
        RECT  4.890 -0.140 5.050 0.660 ;
        RECT  0.700 -0.140 0.980 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.110 0.840 ;
        RECT  0.950 0.680 1.110 1.280 ;
        RECT  2.340 0.660 2.540 1.280 ;
        RECT  0.950 1.120 3.540 1.280 ;
        RECT  0.140 0.300 0.340 1.950 ;
        RECT  3.020 0.300 4.730 0.460 ;
        RECT  3.020 0.300 3.340 0.540 ;
        RECT  4.570 0.300 4.730 1.240 ;
        RECT  4.570 0.960 4.950 1.240 ;
        RECT  3.750 1.080 4.950 1.240 ;
        RECT  3.750 1.080 3.910 1.600 ;
        RECT  3.360 1.440 3.910 1.600 ;
        RECT  1.300 1.760 3.530 1.920 ;
        RECT  3.360 1.440 3.530 2.020 ;
        RECT  3.050 1.760 3.530 2.020 ;
        RECT  5.210 0.360 6.200 0.560 ;
        RECT  6.040 0.360 6.200 1.300 ;
        RECT  5.210 0.360 5.370 1.700 ;
        RECT  4.070 1.540 5.370 1.700 ;
        RECT  4.870 1.540 5.230 2.080 ;
        RECT  4.070 1.540 4.230 2.100 ;
        RECT  3.830 1.940 4.230 2.100 ;
        RECT  6.360 0.410 6.520 1.920 ;
        RECT  5.990 1.640 6.520 1.920 ;
        RECT  8.020 0.920 8.180 1.920 ;
        RECT  5.990 1.760 8.180 1.920 ;
        LAYER VTPH ;
        RECT  6.870 1.080 7.600 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.080 ;
        RECT  0.000 0.000 6.870 1.140 ;
        RECT  7.600 0.000 8.800 1.140 ;
    END
END LACRSM1HM

MACRO LACRSM0HM
    CLASS CORE ;
    FOREIGN LACRSM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.388  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.760 1.900 0.960 ;
        LAYER ME2 ;
        RECT  1.700 0.440 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.320 0.660 2.060 0.960 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        ANTENNAGATEAREA 0.104  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 15.640  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.560 1.240 0.760 1.440 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.760 1.610 ;
        LAYER ME1 ;
        RECT  0.500 1.440 3.060 1.600 ;
        RECT  0.500 1.020 0.790 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.420 0.390 8.700 1.890 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.295  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.240 1.240 7.660 1.600 ;
        RECT  7.460 0.470 7.660 1.600 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 26.880  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.700 0.700 4.410 0.920 ;
        RECT  4.190 0.620 4.410 0.920 ;
        RECT  2.700 0.300 2.860 0.920 ;
        RECT  1.140 0.300 2.860 0.500 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        ANTENNAGATEAREA 0.053  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 10.045  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.580 1.290 5.780 1.490 ;
        LAYER ME2 ;
        RECT  5.300 1.230 5.900 1.570 ;
        LAYER ME1 ;
        RECT  5.530 0.960 5.830 1.680 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  7.860 2.080 8.140 2.540 ;
        RECT  6.780 2.080 7.060 2.540 ;
        RECT  5.590 1.880 5.870 2.540 ;
        RECT  4.390 1.880 4.670 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        RECT  0.740 2.080 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.900 -0.140 8.180 0.660 ;
        RECT  6.900 -0.140 7.180 0.720 ;
        RECT  4.890 -0.140 5.050 0.600 ;
        RECT  0.700 -0.140 0.980 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.110 0.840 ;
        RECT  2.340 0.660 2.540 1.280 ;
        RECT  0.950 0.680 1.110 1.280 ;
        RECT  2.340 1.080 3.540 1.280 ;
        RECT  0.950 1.120 3.540 1.280 ;
        RECT  0.140 0.300 0.340 1.920 ;
        RECT  3.020 0.300 4.730 0.460 ;
        RECT  3.020 0.300 3.300 0.540 ;
        RECT  4.570 0.300 4.730 1.240 ;
        RECT  4.570 0.960 4.950 1.240 ;
        RECT  3.750 1.080 4.950 1.240 ;
        RECT  3.750 1.080 3.910 1.600 ;
        RECT  3.360 1.440 3.910 1.600 ;
        RECT  1.300 1.760 3.530 1.920 ;
        RECT  3.360 1.440 3.530 2.020 ;
        RECT  3.050 1.760 3.530 2.020 ;
        RECT  5.210 0.360 6.200 0.560 ;
        RECT  6.040 0.360 6.200 1.300 ;
        RECT  4.070 1.540 5.370 1.700 ;
        RECT  5.210 0.360 5.370 2.080 ;
        RECT  4.990 1.540 5.370 2.080 ;
        RECT  4.070 1.540 4.230 2.100 ;
        RECT  3.830 1.940 4.230 2.100 ;
        RECT  6.360 0.450 6.520 1.920 ;
        RECT  6.220 1.640 6.520 1.920 ;
        RECT  8.100 0.920 8.260 1.920 ;
        RECT  6.220 1.760 8.260 1.920 ;
        LAYER VTPH ;
        RECT  6.950 1.080 7.860 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.080 ;
        RECT  0.000 0.000 6.950 1.140 ;
        RECT  7.860 0.000 8.800 1.140 ;
    END
END LACRSM0HM

MACRO LACQRSM4HM
    CLASS CORE ;
    FOREIGN LACQRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        ANTENNAGATEAREA 0.092  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 21.835  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.620 0.700 4.240 0.920 ;
        RECT  4.020 0.620 4.240 0.920 ;
        RECT  2.620 0.300 2.780 0.920 ;
        RECT  1.060 0.300 2.780 0.500 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.090  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 0.760 1.500 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.440 1.500 1.160 ;
        LAYER ME1 ;
        RECT  1.240 0.660 1.980 0.960 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.204  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 3.010 1.600 ;
        RECT  0.500 1.020 0.710 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.578  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.840 1.440 7.400 2.070 ;
        RECT  7.200 0.400 7.400 2.070 ;
        RECT  7.010 0.400 7.400 0.690 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        ANTENNAGATEAREA 0.143  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.132  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.420 1.290 5.620 1.490 ;
        LAYER ME2 ;
        RECT  5.420 1.100 5.900 1.680 ;
        LAYER ME1 ;
        RECT  5.360 1.080 5.620 1.680 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.590 1.400 7.820 2.540 ;
        RECT  6.500 1.420 6.660 2.540 ;
        RECT  5.350 1.900 5.630 2.540 ;
        RECT  4.310 1.900 4.590 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.590 -0.140 7.870 0.660 ;
        RECT  6.500 -0.140 6.780 0.680 ;
        RECT  4.720 -0.140 4.880 0.660 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.030 0.840 ;
        RECT  0.870 0.680 1.030 1.280 ;
        RECT  2.260 0.660 2.460 1.280 ;
        RECT  0.870 1.120 3.460 1.280 ;
        RECT  0.140 0.410 0.340 2.080 ;
        RECT  2.940 0.300 4.560 0.460 ;
        RECT  2.940 0.300 3.220 0.540 ;
        RECT  4.400 0.300 4.560 1.240 ;
        RECT  4.400 0.960 4.870 1.240 ;
        RECT  3.620 1.080 4.870 1.240 ;
        RECT  3.620 1.080 3.780 1.600 ;
        RECT  3.280 1.440 3.780 1.600 ;
        RECT  1.220 1.760 3.450 1.920 ;
        RECT  3.280 1.440 3.450 2.020 ;
        RECT  2.970 1.760 3.450 2.020 ;
        RECT  5.040 0.430 5.730 0.630 ;
        RECT  5.540 0.430 5.730 0.920 ;
        RECT  5.540 0.760 6.020 0.920 ;
        RECT  5.830 0.760 6.020 1.300 ;
        RECT  5.040 0.430 5.200 1.700 ;
        RECT  3.940 1.540 5.200 1.700 ;
        RECT  3.940 1.540 4.100 2.100 ;
        RECT  3.660 1.940 4.100 2.100 ;
        RECT  4.790 1.540 5.150 2.100 ;
        RECT  5.930 0.300 6.340 0.600 ;
        RECT  6.180 0.980 7.000 1.260 ;
        RECT  6.180 0.300 6.340 2.100 ;
        RECT  5.870 1.460 6.340 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END LACQRSM4HM

MACRO LACQRSM2HM
    CLASS CORE ;
    FOREIGN LACQRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.090  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 0.760 1.500 0.960 ;
        LAYER ME2 ;
        RECT  1.300 0.440 1.500 1.160 ;
        LAYER ME1 ;
        RECT  1.240 0.660 1.980 0.960 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.092  LAYER ME1  ;
        ANTENNAGATEAREA 0.092  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 22.342  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.620 0.700 4.330 0.920 ;
        RECT  4.070 0.620 4.330 0.920 ;
        RECT  2.620 0.300 2.780 0.920 ;
        RECT  1.060 0.300 2.780 0.500 ;
        END
    END RB
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 3.010 1.600 ;
        RECT  0.500 1.020 0.710 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.449  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.840 1.610 7.500 1.970 ;
        RECT  7.240 0.400 7.500 1.970 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.143  LAYER ME1  ;
        ANTENNAGATEAREA 0.143  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.277  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.510 1.290 5.710 1.490 ;
        LAYER ME2 ;
        RECT  5.300 1.230 5.900 1.570 ;
        LAYER ME1 ;
        RECT  5.450 1.080 5.750 1.680 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.430 2.080 6.710 2.540 ;
        RECT  5.350 1.900 5.630 2.540 ;
        RECT  4.310 1.900 4.590 2.540 ;
        RECT  1.820 2.080 2.100 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.700 -0.140 6.980 0.720 ;
        RECT  4.810 -0.140 4.970 0.660 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.030 0.840 ;
        RECT  0.870 0.680 1.030 1.280 ;
        RECT  2.260 0.660 2.460 1.280 ;
        RECT  0.870 1.120 3.460 1.280 ;
        RECT  0.140 0.300 0.340 1.950 ;
        RECT  2.940 0.300 4.650 0.460 ;
        RECT  2.940 0.300 3.260 0.540 ;
        RECT  4.490 0.300 4.650 1.240 ;
        RECT  4.490 0.960 4.870 1.240 ;
        RECT  3.670 1.080 4.870 1.240 ;
        RECT  3.670 1.080 3.830 1.600 ;
        RECT  3.280 1.440 3.830 1.600 ;
        RECT  1.220 1.760 3.450 1.920 ;
        RECT  3.280 1.440 3.450 2.020 ;
        RECT  2.970 1.760 3.450 2.020 ;
        RECT  5.130 0.430 5.810 0.630 ;
        RECT  5.650 0.430 5.810 0.920 ;
        RECT  5.650 0.760 6.120 0.920 ;
        RECT  5.960 0.760 6.120 1.300 ;
        RECT  5.130 0.430 5.290 1.700 ;
        RECT  3.990 1.540 5.290 1.700 ;
        RECT  3.990 1.540 4.150 2.100 ;
        RECT  3.750 1.940 4.150 2.100 ;
        RECT  4.830 1.540 5.110 2.100 ;
        RECT  6.130 0.300 6.440 0.570 ;
        RECT  6.280 1.060 7.060 1.340 ;
        RECT  6.280 0.300 6.440 1.920 ;
        RECT  5.910 1.640 6.440 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END LACQRSM2HM

MACRO LACQRSM1HM
    CLASS CORE ;
    FOREIGN LACQRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.388  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.760 1.900 0.960 ;
        LAYER ME2 ;
        RECT  1.700 0.440 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.320 0.660 2.060 0.960 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        ANTENNAGATEAREA 0.104  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 15.241  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.590 1.260 0.790 1.460 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.790 1.680 ;
        LAYER ME1 ;
        RECT  0.580 1.440 3.060 1.600 ;
        RECT  0.580 1.020 0.790 1.600 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.150 0.550 7.500 2.040 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.440 1.220 5.900 1.560 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 26.271  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.700 0.700 4.320 0.920 ;
        RECT  4.060 0.620 4.320 0.920 ;
        RECT  2.700 0.300 2.860 0.920 ;
        RECT  1.140 0.300 2.860 0.500 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.690 1.690 6.850 2.540 ;
        RECT  5.520 1.790 5.800 2.540 ;
        RECT  4.360 1.720 4.520 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        RECT  0.740 1.760 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.690 -0.140 6.900 0.860 ;
        RECT  4.800 -0.140 4.960 0.660 ;
        RECT  0.700 -0.140 0.980 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.110 0.840 ;
        RECT  0.950 0.680 1.110 1.280 ;
        RECT  2.340 0.660 2.540 1.280 ;
        RECT  0.950 1.120 3.540 1.280 ;
        RECT  0.140 0.300 0.340 1.950 ;
        RECT  3.020 0.300 4.640 0.460 ;
        RECT  3.020 0.300 3.340 0.540 ;
        RECT  4.480 0.300 4.640 1.240 ;
        RECT  4.480 0.960 4.860 1.240 ;
        RECT  3.700 1.080 4.860 1.240 ;
        RECT  3.700 1.080 3.860 1.600 ;
        RECT  3.360 1.440 3.860 1.600 ;
        RECT  1.300 1.760 3.530 1.920 ;
        RECT  3.360 1.440 3.530 2.020 ;
        RECT  3.050 1.760 3.530 2.020 ;
        RECT  5.120 0.300 6.480 0.460 ;
        RECT  5.580 0.300 5.860 0.640 ;
        RECT  4.020 1.400 5.280 1.560 ;
        RECT  5.120 0.300 5.280 2.010 ;
        RECT  4.880 1.400 5.280 2.010 ;
        RECT  4.020 1.400 4.180 2.100 ;
        RECT  3.740 1.940 4.180 2.100 ;
        RECT  6.060 1.100 6.960 1.380 ;
        RECT  6.060 0.670 6.290 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.520 2.400 ;
        RECT  7.180 1.140 7.600 2.400 ;
        RECT  0.000 1.300 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
        RECT  5.520 0.000 7.180 1.300 ;
    END
END LACQRSM1HM

MACRO LACQRSM0HM
    CLASS CORE ;
    FOREIGN LACQRSM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        ANTENNAGATEAREA 0.104  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 15.241  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.590 1.260 0.790 1.460 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.790 1.680 ;
        LAYER ME1 ;
        RECT  0.580 1.440 3.060 1.600 ;
        RECT  0.580 1.020 0.790 1.600 ;
        END
    END GB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.073  LAYER ME1  ;
        ANTENNAGATEAREA 0.073  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.388  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.760 1.900 0.960 ;
        LAYER ME2 ;
        RECT  1.700 0.440 1.900 1.160 ;
        LAYER ME1 ;
        RECT  1.320 0.660 2.060 0.960 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.150 0.550 7.500 2.040 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.440 1.220 5.900 1.560 ;
        END
    END SB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 26.271  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 0.700 3.900 0.900 ;
        LAYER ME2 ;
        RECT  3.700 0.440 3.900 1.160 ;
        LAYER ME1 ;
        RECT  2.700 0.700 4.320 0.920 ;
        RECT  4.060 0.620 4.320 0.920 ;
        RECT  2.700 0.300 2.860 0.920 ;
        RECT  1.140 0.300 2.860 0.500 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.660 1.690 6.820 2.540 ;
        RECT  5.520 1.790 5.800 2.540 ;
        RECT  4.360 1.720 4.520 2.540 ;
        RECT  1.900 2.080 2.180 2.540 ;
        RECT  0.740 1.760 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.660 -0.140 6.870 0.860 ;
        RECT  4.800 -0.140 4.960 0.660 ;
        RECT  0.700 -0.140 0.980 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.680 1.110 0.840 ;
        RECT  0.950 0.680 1.110 1.280 ;
        RECT  2.340 0.660 2.540 1.280 ;
        RECT  0.950 1.120 3.540 1.280 ;
        RECT  0.140 0.300 0.340 1.950 ;
        RECT  3.020 0.300 4.640 0.460 ;
        RECT  3.020 0.300 3.340 0.540 ;
        RECT  4.480 0.300 4.640 1.240 ;
        RECT  4.480 0.960 4.860 1.240 ;
        RECT  3.700 1.080 4.860 1.240 ;
        RECT  3.700 1.080 3.860 1.600 ;
        RECT  3.360 1.440 3.860 1.600 ;
        RECT  1.300 1.760 3.530 1.920 ;
        RECT  3.360 1.440 3.530 2.020 ;
        RECT  3.050 1.760 3.530 2.020 ;
        RECT  5.120 0.300 6.430 0.460 ;
        RECT  4.020 1.400 5.280 1.560 ;
        RECT  5.120 0.300 5.280 2.010 ;
        RECT  4.880 1.400 5.280 2.010 ;
        RECT  4.020 1.400 4.180 2.100 ;
        RECT  3.740 1.940 4.180 2.100 ;
        RECT  6.060 1.100 6.930 1.380 ;
        RECT  6.060 0.670 6.280 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.520 2.400 ;
        RECT  7.140 1.140 7.600 2.400 ;
        RECT  0.000 1.300 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
        RECT  5.520 0.000 7.140 1.300 ;
    END
END LACQRSM0HM

MACRO LACQM4HM
    CLASS CORE ;
    FOREIGN LACQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.400 0.420 5.720 2.100 ;
        RECT  5.240 0.840 5.720 1.160 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  6.000 1.410 6.200 2.540 ;
        RECT  4.960 1.410 5.160 2.540 ;
        RECT  3.700 1.820 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.980 -0.140 6.180 0.680 ;
        RECT  4.940 -0.140 5.140 0.680 ;
        RECT  3.940 -0.140 4.140 0.580 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  3.480 1.060 3.640 1.660 ;
        RECT  4.480 0.380 4.640 1.660 ;
        RECT  3.480 1.500 4.640 1.660 ;
        RECT  4.170 1.500 4.460 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END LACQM4HM

MACRO LACQM2HM
    CLASS CORE ;
    FOREIGN LACQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.420 5.160 1.910 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.480 1.640 5.680 2.540 ;
        RECT  3.660 1.810 3.940 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.460 -0.140 5.660 0.680 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  4.380 0.340 4.740 0.500 ;
        RECT  3.480 1.060 3.640 1.650 ;
        RECT  3.480 1.490 4.540 1.650 ;
        RECT  4.380 0.340 4.540 2.100 ;
        RECT  4.240 1.490 4.540 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END LACQM2HM

MACRO LACQM1HM
    CLASS CORE ;
    FOREIGN LACQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.460 5.160 1.780 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.480 1.640 5.680 2.540 ;
        RECT  3.660 1.810 3.940 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.460 -0.140 5.660 0.680 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  4.380 0.340 4.740 0.500 ;
        RECT  3.480 1.060 3.640 1.650 ;
        RECT  3.480 1.490 4.540 1.650 ;
        RECT  4.380 0.340 4.540 2.100 ;
        RECT  4.240 1.490 4.540 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END LACQM1HM

MACRO LACQM0HM
    CLASS CORE ;
    FOREIGN LACQM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.245  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 0.470 5.160 1.780 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.480 1.640 5.680 2.540 ;
        RECT  3.660 1.810 3.940 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.420 -0.140 5.700 0.680 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  4.380 0.340 4.740 0.500 ;
        RECT  3.480 1.060 3.640 1.650 ;
        RECT  3.480 1.490 4.540 1.650 ;
        RECT  4.380 0.340 4.540 2.100 ;
        RECT  4.240 1.490 4.540 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END LACQM0HM

MACRO LACM4HM
    CLASS CORE ;
    FOREIGN LACM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.550  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.220 0.900 5.660 1.100 ;
        RECT  5.460 0.420 5.660 1.100 ;
        RECT  5.220 0.900 5.380 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.380 1.400 6.780 1.600 ;
        RECT  6.620 0.400 6.780 1.600 ;
        RECT  6.500 0.400 6.780 0.760 ;
        RECT  6.380 1.400 6.580 2.100 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.880 1.760 7.080 2.540 ;
        RECT  5.860 1.640 6.060 2.540 ;
        RECT  4.540 1.920 4.740 2.540 ;
        RECT  3.700 1.820 3.900 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.020 -0.140 7.220 0.680 ;
        RECT  5.980 -0.140 6.180 0.680 ;
        RECT  4.940 -0.140 5.140 0.680 ;
        RECT  3.940 -0.140 4.140 0.580 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.320 0.900 ;
        RECT  4.160 0.740 4.320 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  6.060 1.060 6.460 1.220 ;
        RECT  6.060 1.060 6.220 1.480 ;
        RECT  5.540 1.320 6.220 1.480 ;
        RECT  3.480 1.060 3.640 1.660 ;
        RECT  4.480 0.380 4.640 1.660 ;
        RECT  3.480 1.500 5.060 1.660 ;
        RECT  4.900 1.500 5.060 2.100 ;
        RECT  5.540 1.320 5.700 2.100 ;
        RECT  4.900 1.940 5.700 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END LACM4HM

MACRO LACM2HM
    CLASS CORE ;
    FOREIGN LACM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.503  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.960 0.420 5.160 1.100 ;
        RECT  4.840 0.900 5.000 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.000 0.400 6.300 2.100 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.480 1.640 5.680 2.540 ;
        RECT  3.660 1.810 3.940 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.460 -0.140 5.660 0.680 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  4.380 0.340 4.740 0.500 ;
        RECT  5.660 0.960 5.820 1.480 ;
        RECT  5.160 1.320 5.820 1.480 ;
        RECT  3.480 1.060 3.640 1.650 ;
        RECT  3.480 1.490 4.540 1.650 ;
        RECT  4.380 0.340 4.540 2.100 ;
        RECT  4.240 1.490 4.540 2.100 ;
        RECT  5.160 1.320 5.320 2.100 ;
        RECT  4.240 1.940 5.320 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END LACM2HM

MACRO LACM1HM
    CLASS CORE ;
    FOREIGN LACM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.353  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.960 0.460 5.160 1.100 ;
        RECT  4.840 0.900 5.000 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.000 0.440 6.300 1.820 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.480 1.640 5.680 2.540 ;
        RECT  3.660 1.810 3.940 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.460 -0.140 5.660 0.680 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  4.380 0.340 4.740 0.500 ;
        RECT  5.660 0.960 5.820 1.480 ;
        RECT  5.160 1.320 5.820 1.480 ;
        RECT  3.480 1.060 3.640 1.650 ;
        RECT  3.480 1.490 4.540 1.650 ;
        RECT  4.380 0.340 4.540 2.100 ;
        RECT  4.240 1.490 4.540 2.100 ;
        RECT  5.160 1.320 5.320 2.100 ;
        RECT  4.240 1.940 5.320 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END LACM1HM

MACRO LACM0HM
    CLASS CORE ;
    FOREIGN LACM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 0.840 2.300 1.160 ;
        END
    END D
    PIN GB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END GB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.295  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.960 0.470 5.160 1.100 ;
        RECT  4.800 0.900 5.000 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.245  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.000 0.440 6.300 1.850 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.480 1.640 5.680 2.540 ;
        RECT  3.660 1.810 3.940 2.540 ;
        RECT  1.700 1.640 1.980 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.420 -0.140 5.700 0.680 ;
        RECT  3.940 -0.140 4.140 0.560 ;
        RECT  1.740 -0.140 1.940 0.560 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.100 0.680 ;
        RECT  0.940 0.520 1.100 1.480 ;
        RECT  0.160 1.320 1.100 1.480 ;
        RECT  0.160 1.320 0.320 1.840 ;
        RECT  3.100 0.620 3.420 0.900 ;
        RECT  1.280 1.320 2.620 1.480 ;
        RECT  1.280 0.320 1.440 1.840 ;
        RECT  2.460 1.020 2.620 2.100 ;
        RECT  3.100 0.620 3.260 2.100 ;
        RECT  2.460 1.940 3.260 2.100 ;
        RECT  2.580 0.300 3.740 0.460 ;
        RECT  2.580 0.300 2.940 0.520 ;
        RECT  3.580 0.300 3.740 0.900 ;
        RECT  3.580 0.740 4.220 0.900 ;
        RECT  4.060 0.740 4.220 1.320 ;
        RECT  2.780 0.300 2.940 1.760 ;
        RECT  4.380 0.340 4.740 0.500 ;
        RECT  5.660 0.960 5.820 1.480 ;
        RECT  5.160 1.320 5.820 1.480 ;
        RECT  3.480 1.060 3.640 1.650 ;
        RECT  3.480 1.490 4.540 1.650 ;
        RECT  4.380 0.340 4.540 2.100 ;
        RECT  4.240 1.490 4.540 2.100 ;
        RECT  5.160 1.320 5.320 2.100 ;
        RECT  4.240 1.940 5.320 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END LACM0HM

MACRO INVM8HM
    CLASS CORE ;
    FOREIGN INVM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.500 1.320 ;
        RECT  0.100 0.840 0.360 1.320 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.410 1.900 1.970 ;
        RECT  0.620 1.520 1.900 1.720 ;
        RECT  1.660 0.680 1.900 1.720 ;
        RECT  0.660 0.680 1.900 0.880 ;
        RECT  0.620 1.520 0.860 2.000 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.610 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END INVM8HM

MACRO INVM6HM
    CLASS CORE ;
    FOREIGN INVM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.500 1.320 ;
        RECT  0.100 0.840 0.360 1.320 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.410 1.900 1.880 ;
        RECT  0.660 1.540 1.900 1.740 ;
        RECT  0.660 0.680 1.900 0.880 ;
        RECT  0.660 1.540 0.860 1.910 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END INVM6HM

MACRO INVM5HM
    CLASS CORE ;
    FOREIGN INVM5HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.500 1.320 ;
        RECT  0.100 0.840 0.360 1.320 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.770  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.410 1.900 1.960 ;
        RECT  0.620 1.540 1.900 1.740 ;
        RECT  0.660 0.680 1.900 0.880 ;
        RECT  0.620 1.540 0.860 1.990 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.720 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END INVM5HM

MACRO INVM4HM
    CLASS CORE ;
    FOREIGN INVM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.050 1.100 1.320 ;
        RECT  0.100 0.840 0.360 1.320 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.620 1.480 1.500 1.680 ;
        RECT  1.300 0.680 1.500 1.680 ;
        RECT  0.660 0.680 1.500 0.880 ;
        RECT  0.620 1.480 0.900 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END INVM4HM

MACRO INVM48HM
    CLASS CORE ;
    FOREIGN INVM48HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 6.037  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.422  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.764  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.990 5.900 1.270 ;
        RECT  0.100 0.990 0.400 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.878  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.060 1.480 12.340 2.100 ;
        RECT  0.620 0.670 12.340 0.830 ;
        RECT  12.060 0.310 12.340 0.830 ;
        RECT  0.620 1.480 12.340 1.740 ;
        RECT  11.020 1.480 11.300 2.100 ;
        RECT  11.020 0.300 11.300 0.830 ;
        RECT  9.980 1.480 10.260 2.100 ;
        RECT  9.980 0.390 10.260 0.830 ;
        RECT  8.940 1.480 9.220 2.100 ;
        RECT  8.940 0.390 9.220 0.830 ;
        RECT  7.900 1.480 8.180 2.100 ;
        RECT  7.900 0.390 8.180 0.830 ;
        RECT  6.860 1.480 7.140 2.100 ;
        RECT  0.620 0.660 7.140 0.830 ;
        RECT  6.860 0.390 7.140 0.830 ;
        RECT  6.110 0.660 6.710 1.740 ;
        RECT  5.820 1.480 6.100 2.100 ;
        RECT  5.820 0.390 6.100 0.830 ;
        RECT  4.780 1.480 5.060 2.100 ;
        RECT  4.780 0.390 5.060 0.830 ;
        RECT  3.740 1.480 4.020 2.100 ;
        RECT  3.740 0.390 4.020 0.830 ;
        RECT  2.700 1.480 2.980 2.100 ;
        RECT  2.700 0.390 2.980 0.830 ;
        RECT  1.660 1.480 1.940 2.100 ;
        RECT  1.660 0.390 1.940 0.830 ;
        RECT  0.620 1.480 0.900 2.100 ;
        RECT  0.620 0.390 0.900 0.830 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.540 1.900 11.820 2.540 ;
        RECT  10.500 1.900 10.780 2.540 ;
        RECT  9.460 1.900 9.740 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.880 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.540 -0.140 11.820 0.500 ;
        RECT  10.500 -0.140 10.780 0.500 ;
        RECT  9.460 -0.140 9.740 0.500 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.100 -0.140 0.380 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  6.900 0.990 11.860 1.270 ;
        LAYER VTPH ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
    END
END INVM48HM

MACRO INVM40HM
    CLASS CORE ;
    FOREIGN INVM40HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 4.774  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.827  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.688  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 5.100 1.300 ;
        RECT  0.100 0.840 0.360 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.886  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.020 1.460 10.260 2.100 ;
        RECT  0.660 0.660 10.220 0.860 ;
        RECT  10.020 0.300 10.220 0.860 ;
        RECT  0.620 1.460 10.260 1.720 ;
        RECT  8.980 1.460 9.180 2.100 ;
        RECT  8.980 0.390 9.180 0.860 ;
        RECT  7.940 1.460 8.140 2.100 ;
        RECT  7.940 0.390 8.140 0.860 ;
        RECT  6.900 1.460 7.100 2.100 ;
        RECT  6.900 0.390 7.100 0.860 ;
        RECT  5.860 1.460 6.060 2.100 ;
        RECT  5.860 0.390 6.060 0.860 ;
        RECT  5.300 0.660 5.900 1.720 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.390 5.020 0.860 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.390 3.980 0.860 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.390 2.940 0.860 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.390 1.900 0.860 ;
        RECT  0.620 1.460 0.860 2.100 ;
        RECT  0.660 0.390 0.860 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.460 1.880 9.740 2.540 ;
        RECT  8.420 1.880 8.700 2.540 ;
        RECT  7.380 1.880 7.660 2.540 ;
        RECT  6.340 1.880 6.620 2.540 ;
        RECT  5.300 1.880 5.580 2.540 ;
        RECT  4.260 1.880 4.540 2.540 ;
        RECT  3.220 1.880 3.500 2.540 ;
        RECT  2.180 1.880 2.460 2.540 ;
        RECT  1.140 1.880 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.460 -0.140 9.740 0.500 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  6.100 1.080 9.620 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.140 ;
    END
END INVM40HM

MACRO INVM3HM
    CLASS CORE ;
    FOREIGN INVM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.223  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.100 1.320 ;
        RECT  0.100 0.840 0.360 1.320 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.372  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.510 1.500 1.710 ;
        RECT  1.300 0.680 1.500 1.710 ;
        RECT  0.660 0.680 1.500 0.880 ;
        RECT  0.660 1.510 0.860 2.050 ;
        RECT  0.660 0.350 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.140 1.870 1.420 2.540 ;
        RECT  0.140 1.780 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END INVM3HM

MACRO INVM36HM
    CLASS CORE ;
    FOREIGN INVM36HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 4.472  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.678  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.670  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.090 1.080 4.510 1.300 ;
        RECT  0.090 0.840 0.400 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.464  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.980 1.460 9.220 2.100 ;
        RECT  0.660 0.680 9.180 0.880 ;
        RECT  8.980 0.430 9.180 0.880 ;
        RECT  0.620 1.460 9.220 1.740 ;
        RECT  7.940 1.460 8.140 2.100 ;
        RECT  7.940 0.430 8.140 0.880 ;
        RECT  6.900 1.460 7.100 2.100 ;
        RECT  6.900 0.430 7.100 0.880 ;
        RECT  5.860 1.460 6.060 2.100 ;
        RECT  5.860 0.430 6.060 0.880 ;
        RECT  4.900 0.680 5.500 1.740 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.430 5.020 0.880 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.430 3.980 0.880 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.430 2.940 0.880 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.430 1.900 0.880 ;
        RECT  0.620 1.460 0.860 2.100 ;
        RECT  0.660 0.430 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.460 1.460 9.740 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.460 -0.140 9.740 0.630 ;
        RECT  8.420 -0.140 8.700 0.520 ;
        RECT  7.380 -0.140 7.660 0.520 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  5.700 1.080 9.220 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
    END
END INVM36HM

MACRO INVM32HM
    CLASS CORE ;
    FOREIGN INVM32HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 3.962  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.381  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.664  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 3.900 1.300 ;
        RECT  0.100 0.840 0.400 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.968  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.940 1.460 8.180 2.100 ;
        RECT  0.660 0.680 8.140 0.880 ;
        RECT  7.940 0.410 8.140 0.880 ;
        RECT  0.620 1.460 8.180 1.720 ;
        RECT  6.900 1.460 7.100 2.100 ;
        RECT  6.900 0.410 7.100 0.880 ;
        RECT  5.860 1.460 6.060 2.100 ;
        RECT  5.860 0.410 6.060 0.880 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  4.100 0.680 4.700 1.720 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.410 3.980 0.880 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.410 2.940 0.880 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  0.620 1.460 0.860 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.420 1.880 8.700 2.540 ;
        RECT  7.380 1.880 7.660 2.540 ;
        RECT  6.340 1.880 6.620 2.540 ;
        RECT  5.300 1.880 5.580 2.540 ;
        RECT  4.260 1.880 4.540 2.540 ;
        RECT  3.220 1.880 3.500 2.540 ;
        RECT  2.180 1.880 2.460 2.540 ;
        RECT  1.140 1.880 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.420 -0.140 8.700 0.520 ;
        RECT  7.380 -0.140 7.660 0.520 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.900 1.080 8.060 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END INVM32HM

MACRO INVM2HM
    CLASS CORE ;
    FOREIGN INVM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.450 1.100 2.090 ;
        RECT  0.900 0.370 1.100 2.090 ;
        RECT  0.720 0.370 1.100 0.570 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.270 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.200 1.480 0.480 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.240 -0.140 0.440 0.610 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END INVM2HM

MACRO INVM28HM
    CLASS CORE ;
    FOREIGN INVM28HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 3.557  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.083  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.707  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 3.500 1.280 ;
        RECT  0.100 0.840 0.400 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.900 1.460 7.140 2.100 ;
        RECT  0.660 0.680 7.100 0.880 ;
        RECT  6.900 0.410 7.100 0.880 ;
        RECT  0.620 1.460 7.140 1.740 ;
        RECT  5.860 1.460 6.060 2.100 ;
        RECT  5.860 0.410 6.060 0.880 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  3.700 0.680 4.300 1.740 ;
        RECT  3.780 0.410 3.980 2.100 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.410 2.940 0.880 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  0.620 1.460 0.860 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.560 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.380 -0.140 7.660 0.520 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.500 1.080 7.300 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END INVM28HM

MACRO INVM24HM
    CLASS CORE ;
    FOREIGN INVM24HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.974  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.786  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.666  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 3.100 1.280 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.976  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.820 1.460 6.100 2.100 ;
        RECT  0.660 0.680 6.060 0.880 ;
        RECT  5.860 0.410 6.060 0.880 ;
        RECT  0.620 1.460 6.100 1.740 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.410 3.980 0.880 ;
        RECT  0.620 1.440 3.900 1.740 ;
        RECT  3.300 0.680 3.900 1.740 ;
        RECT  2.740 1.440 2.940 2.100 ;
        RECT  2.740 0.410 2.940 0.880 ;
        RECT  1.700 1.440 1.900 2.100 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  0.620 1.440 0.860 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.520 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.100 1.080 6.180 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END INVM24HM

MACRO INVM20HM
    CLASS CORE ;
    FOREIGN INVM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.402  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.488  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.615  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 2.700 1.300 ;
        RECT  0.100 0.840 0.500 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.480  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.460 5.060 2.100 ;
        RECT  0.660 0.680 5.020 0.880 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  0.620 1.460 5.060 1.740 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.410 3.980 0.880 ;
        RECT  2.900 0.680 3.500 1.740 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.410 2.940 0.880 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  0.620 1.460 0.860 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.300 1.500 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.700 1.080 5.060 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END INVM20HM

MACRO INVM1HM
    CLASS CORE ;
    FOREIGN INVM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.560 1.100 1.860 ;
        RECT  0.900 0.400 1.100 1.860 ;
        RECT  0.720 0.400 1.100 0.600 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.400 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.240 1.560 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.240 -0.140 0.440 0.600 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END INVM1HM

MACRO INVM18HM
    CLASS CORE ;
    FOREIGN INVM18HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.205  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.339  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.646  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 2.300 1.320 ;
        RECT  0.100 0.840 0.460 1.320 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.406  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.520 5.060 2.100 ;
        RECT  0.660 0.680 5.020 0.880 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  0.620 1.520 5.060 1.740 ;
        RECT  3.780 1.520 3.980 2.100 ;
        RECT  3.780 0.410 3.980 0.880 ;
        RECT  2.500 0.680 3.100 1.740 ;
        RECT  2.740 0.410 2.940 2.100 ;
        RECT  1.700 1.520 1.900 2.100 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  0.620 1.520 0.860 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.300 1.080 4.660 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END INVM18HM

MACRO INVM16HM
    CLASS CORE ;
    FOREIGN INVM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.815  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.190  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.525  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.900 1.330 ;
        RECT  0.100 0.840 0.400 1.330 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.740 1.540 4.060 2.100 ;
        RECT  0.660 0.680 3.980 0.880 ;
        RECT  3.780 0.410 3.980 0.880 ;
        RECT  0.620 1.540 4.060 1.740 ;
        RECT  2.700 1.540 2.980 2.100 ;
        RECT  2.740 0.410 2.940 0.880 ;
        RECT  2.100 0.680 2.700 1.740 ;
        RECT  1.660 1.540 1.940 2.100 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  0.620 1.540 0.900 2.100 ;
        RECT  0.660 0.410 0.860 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.260 1.510 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.490 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.260 -0.140 4.540 0.660 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.080 3.900 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END INVM16HM

MACRO INVM14HM
    CLASS CORE ;
    FOREIGN INVM14HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.591  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.042  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.528  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 1.500 1.300 ;
        RECT  0.100 0.840 0.310 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.910  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.500 4.020 2.080 ;
        RECT  0.660 0.660 3.980 0.840 ;
        RECT  3.780 0.390 3.980 0.840 ;
        RECT  0.620 1.500 4.020 1.700 ;
        RECT  2.740 1.500 2.940 2.080 ;
        RECT  2.740 0.390 2.940 0.840 ;
        RECT  1.700 0.660 2.300 1.700 ;
        RECT  1.700 0.390 1.900 2.080 ;
        RECT  0.620 1.500 0.860 2.080 ;
        RECT  0.660 0.390 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.500 1.040 3.500 1.240 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END INVM14HM

MACRO INVM12HM
    CLASS CORE ;
    FOREIGN INVM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.446  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.619  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 1.500 1.300 ;
        RECT  0.100 0.840 0.300 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.500 2.980 2.080 ;
        RECT  0.660 0.660 2.940 0.840 ;
        RECT  2.740 0.390 2.940 0.840 ;
        RECT  0.620 1.500 2.980 1.700 ;
        RECT  1.700 0.660 2.300 1.700 ;
        RECT  1.700 0.390 1.900 2.080 ;
        RECT  0.620 1.500 0.860 2.080 ;
        RECT  0.660 0.390 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.500 1.000 3.140 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END INVM12HM

MACRO INVM10HM
    CLASS CORE ;
    FOREIGN INVM10HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.420  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.744  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.908  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 1.450 1.300 ;
        RECT  0.100 0.840 0.300 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.414  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 1.500 3.080 2.080 ;
        RECT  0.760 0.660 3.040 0.840 ;
        RECT  2.840 0.390 3.040 0.840 ;
        RECT  0.720 1.500 3.080 1.700 ;
        RECT  1.800 1.500 2.000 2.080 ;
        RECT  1.800 0.390 2.000 0.840 ;
        RECT  1.640 0.660 1.960 1.700 ;
        RECT  0.720 1.500 0.960 2.080 ;
        RECT  0.760 0.390 0.960 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.280 1.900 2.560 2.540 ;
        RECT  1.240 1.900 1.520 2.540 ;
        RECT  0.200 1.500 0.480 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.280 -0.140 2.560 0.500 ;
        RECT  1.240 -0.140 1.520 0.500 ;
        RECT  0.240 -0.140 0.440 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.120 1.000 2.740 1.300 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END INVM10HM

MACRO INVM0HM
    CLASS CORE ;
    FOREIGN INVM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.520 1.100 1.820 ;
        RECT  0.900 0.440 1.100 1.820 ;
        RECT  0.720 0.440 1.100 0.640 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.360 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.240 1.520 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.240 -0.140 0.440 0.680 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END INVM0HM

MACRO FILE8HM
    CLASS CORE ;
    FOREIGN FILE8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.340 1.730 2.540 2.540 ;
        RECT  0.620 1.660 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.300 -0.140 2.580 0.540 ;
        RECT  0.660 -0.140 0.860 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.180 0.560 1.380 ;
        RECT  0.140 1.180 0.340 1.880 ;
        RECT  0.140 0.340 0.340 0.980 ;
        RECT  0.140 0.780 0.920 0.980 ;
        RECT  0.720 0.780 0.920 1.460 ;
        RECT  0.720 1.260 2.080 1.460 ;
        RECT  1.080 0.740 2.440 0.940 ;
        RECT  2.240 0.740 2.440 1.430 ;
        RECT  2.240 1.230 3.060 1.430 ;
        RECT  2.860 1.230 3.060 2.010 ;
        RECT  2.860 0.300 3.060 0.990 ;
        RECT  2.640 0.790 3.060 0.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END FILE8HM

MACRO FILE64HM
    CLASS CORE ;
    FOREIGN FILE64HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 25.600 2.540 ;
        RECT  24.740 1.730 24.940 2.540 ;
        RECT  21.730 1.730 21.930 2.540 ;
        RECT  18.720 1.730 18.920 2.540 ;
        RECT  15.710 1.730 15.910 2.540 ;
        RECT  12.700 1.730 12.900 2.540 ;
        RECT  9.690 1.730 9.890 2.540 ;
        RECT  6.680 1.730 6.880 2.540 ;
        RECT  3.670 1.730 3.870 2.540 ;
        RECT  0.660 1.600 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 25.600 0.140 ;
        RECT  24.700 -0.140 24.980 0.540 ;
        RECT  21.690 -0.140 21.970 0.540 ;
        RECT  18.680 -0.140 18.960 0.540 ;
        RECT  15.670 -0.140 15.950 0.540 ;
        RECT  12.660 -0.140 12.940 0.540 ;
        RECT  9.650 -0.140 9.930 0.540 ;
        RECT  6.640 -0.140 6.920 0.540 ;
        RECT  3.630 -0.140 3.910 0.540 ;
        RECT  0.660 -0.140 0.860 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.180 0.560 1.380 ;
        RECT  0.140 1.180 0.340 1.880 ;
        RECT  0.140 0.340 0.340 0.980 ;
        RECT  0.140 0.780 1.160 0.980 ;
        RECT  0.960 0.780 1.160 1.460 ;
        RECT  0.960 1.260 24.470 1.460 ;
        RECT  1.320 0.740 24.830 0.940 ;
        RECT  24.630 0.740 24.830 1.430 ;
        RECT  24.630 1.230 25.460 1.430 ;
        RECT  25.260 1.230 25.460 2.010 ;
        RECT  25.260 0.300 25.460 0.990 ;
        RECT  25.040 0.790 25.460 0.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 25.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 25.600 1.140 ;
    END
END FILE64HM

MACRO FILE4HM
    CLASS CORE ;
    FOREIGN FILE4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.260 1.710 1.460 2.540 ;
        RECT  0.660 1.710 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.740 -0.140 0.940 0.590 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.760 1.080 0.960 ;
        RECT  0.140 0.760 0.340 1.980 ;
        RECT  1.260 0.320 1.460 1.440 ;
        RECT  0.520 1.240 1.460 1.440 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END FILE4HM

MACRO FILE3HM
    CLASS CORE ;
    FOREIGN FILE3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.860 1.710 1.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.720 0.700 1.000 ;
        RECT  0.140 0.720 0.340 1.990 ;
        RECT  0.860 0.320 1.060 1.480 ;
        RECT  0.500 1.200 1.060 1.480 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END FILE3HM

MACRO FILE32HM
    CLASS CORE ;
    FOREIGN FILE32HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.940 1.730 12.140 2.540 ;
        RECT  9.120 1.730 9.320 2.540 ;
        RECT  6.300 1.730 6.500 2.540 ;
        RECT  3.480 1.730 3.680 2.540 ;
        RECT  0.660 1.600 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.900 -0.140 12.180 0.540 ;
        RECT  9.080 -0.140 9.360 0.540 ;
        RECT  6.260 -0.140 6.540 0.540 ;
        RECT  3.440 -0.140 3.720 0.540 ;
        RECT  0.660 -0.140 0.860 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.180 0.560 1.380 ;
        RECT  0.140 1.180 0.340 1.880 ;
        RECT  0.140 0.320 0.340 0.980 ;
        RECT  0.140 0.780 1.160 0.980 ;
        RECT  0.960 0.780 1.160 1.460 ;
        RECT  0.960 1.260 11.680 1.460 ;
        RECT  1.320 0.740 12.040 0.940 ;
        RECT  11.840 0.740 12.040 1.430 ;
        RECT  11.840 1.230 12.660 1.430 ;
        RECT  12.460 1.230 12.660 2.010 ;
        RECT  12.460 0.300 12.660 0.990 ;
        RECT  12.240 0.790 12.660 0.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
    END
END FILE32HM

MACRO FILE16HM
    CLASS CORE ;
    FOREIGN FILE16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.540 1.730 5.740 2.540 ;
        RECT  3.100 1.730 3.300 2.540 ;
        RECT  0.660 1.600 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.500 -0.140 5.780 0.540 ;
        RECT  3.060 -0.140 3.340 0.540 ;
        RECT  0.660 -0.140 0.860 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.180 0.560 1.380 ;
        RECT  0.140 1.180 0.340 1.880 ;
        RECT  0.140 0.320 0.340 0.980 ;
        RECT  0.140 0.780 1.160 0.980 ;
        RECT  0.960 0.780 1.160 1.460 ;
        RECT  0.960 1.260 5.280 1.460 ;
        RECT  1.640 0.740 5.640 0.940 ;
        RECT  5.440 0.740 5.640 1.430 ;
        RECT  5.440 1.230 6.260 1.430 ;
        RECT  6.060 1.230 6.260 2.010 ;
        RECT  6.060 0.300 6.260 0.990 ;
        RECT  5.840 0.790 6.260 0.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END FILE16HM

MACRO FILE128HM
    CLASS CORE ;
    FOREIGN FILE128HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 51.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 51.200 2.540 ;
        RECT  50.300 1.730 50.500 2.540 ;
        RECT  47.200 1.730 47.400 2.540 ;
        RECT  44.100 1.730 44.300 2.540 ;
        RECT  41.000 1.730 41.200 2.540 ;
        RECT  37.900 1.730 38.100 2.540 ;
        RECT  34.800 1.730 35.000 2.540 ;
        RECT  31.700 1.730 31.900 2.540 ;
        RECT  28.600 1.730 28.800 2.540 ;
        RECT  25.500 1.730 25.700 2.540 ;
        RECT  22.400 1.730 22.600 2.540 ;
        RECT  19.300 1.730 19.500 2.540 ;
        RECT  16.200 1.730 16.400 2.540 ;
        RECT  13.100 1.730 13.300 2.540 ;
        RECT  10.000 1.730 10.200 2.540 ;
        RECT  6.900 1.730 7.100 2.540 ;
        RECT  3.800 1.730 4.000 2.540 ;
        RECT  0.700 1.600 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 51.200 0.140 ;
        RECT  50.260 -0.140 50.540 0.540 ;
        RECT  47.160 -0.140 47.440 0.540 ;
        RECT  44.060 -0.140 44.350 0.540 ;
        RECT  40.960 -0.140 41.240 0.540 ;
        RECT  37.860 -0.140 38.140 0.540 ;
        RECT  34.760 -0.140 35.040 0.540 ;
        RECT  31.660 -0.140 31.940 0.540 ;
        RECT  28.560 -0.140 28.840 0.540 ;
        RECT  25.460 -0.140 25.740 0.540 ;
        RECT  22.360 -0.140 22.640 0.540 ;
        RECT  19.260 -0.140 19.540 0.540 ;
        RECT  16.160 -0.140 16.440 0.540 ;
        RECT  13.060 -0.140 13.340 0.540 ;
        RECT  9.960 -0.140 10.240 0.540 ;
        RECT  6.860 -0.140 7.140 0.540 ;
        RECT  3.760 -0.140 4.040 0.540 ;
        RECT  0.700 -0.140 0.900 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 1.180 0.600 1.380 ;
        RECT  0.180 1.180 0.380 1.880 ;
        RECT  0.180 0.320 0.380 0.980 ;
        RECT  0.180 0.780 1.250 0.980 ;
        RECT  1.050 0.780 1.250 1.460 ;
        RECT  1.050 1.260 50.070 1.460 ;
        RECT  1.490 0.740 50.440 0.940 ;
        RECT  50.240 0.740 50.440 1.430 ;
        RECT  50.240 1.230 51.020 1.430 ;
        RECT  50.820 1.230 51.020 2.010 ;
        RECT  50.820 0.320 51.020 0.990 ;
        RECT  50.600 0.790 51.020 0.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 51.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 51.200 1.140 ;
    END
END FILE128HM

MACRO FIL8HM
    CLASS CORE ;
    FOREIGN FIL8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END FIL8HM

MACRO FIL64HM
    CLASS CORE ;
    FOREIGN FIL64HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 25.600 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 25.600 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 25.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 25.600 1.140 ;
    END
END FIL64HM

MACRO FIL4HM
    CLASS CORE ;
    FOREIGN FIL4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END FIL4HM

MACRO FIL32HM
    CLASS CORE ;
    FOREIGN FIL32HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
    END
END FIL32HM

MACRO FIL2HM
    CLASS CORE ;
    FOREIGN FIL2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.800 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.800 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.800 1.140 ;
    END
END FIL2HM

MACRO FIL1HM
    CLASS CORE ;
    FOREIGN FIL1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.400 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.400 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.400 1.140 ;
    END
END FIL1HM

MACRO FIL16HM
    CLASS CORE ;
    FOREIGN FIL16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END FIL16HM

MACRO DFZRM8HM
    CLASS CORE ;
    FOREIGN DFZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.265  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.630 0.900 11.350 1.200 ;
        RECT  11.070 0.620 11.350 1.200 ;
        RECT  11.070 0.620 11.230 1.760 ;
        RECT  9.750 0.620 9.910 1.760 ;
        RECT  9.630 0.620 9.910 1.200 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.890 0.440 15.100 2.080 ;
        RECT  13.850 1.440 15.100 1.640 ;
        RECT  13.850 0.720 15.100 0.920 ;
        RECT  13.850 1.440 14.050 2.080 ;
        RECT  13.850 0.440 14.050 0.920 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.000 2.540 ;
        RECT  15.410 1.440 15.610 2.540 ;
        RECT  14.370 1.840 14.570 2.540 ;
        RECT  13.240 1.480 13.440 2.540 ;
        RECT  11.710 1.900 11.990 2.540 ;
        RECT  10.390 1.840 10.590 2.540 ;
        RECT  9.070 1.840 9.270 2.540 ;
        RECT  7.750 2.020 7.950 2.540 ;
        RECT  4.790 2.080 5.070 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.000 0.140 ;
        RECT  15.410 -0.140 15.610 0.720 ;
        RECT  14.370 -0.140 14.570 0.560 ;
        RECT  13.350 -0.140 13.510 0.650 ;
        RECT  11.830 -0.140 12.110 0.320 ;
        RECT  10.390 -0.140 10.590 0.380 ;
        RECT  8.900 -0.140 9.100 0.660 ;
        RECT  7.710 -0.140 7.990 0.320 ;
        RECT  4.790 -0.140 5.070 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.710 0.920 5.330 1.080 ;
        RECT  3.710 0.640 3.990 1.780 ;
        RECT  4.370 1.240 5.750 1.400 ;
        RECT  5.550 0.620 5.750 1.780 ;
        RECT  0.140 0.400 0.340 0.680 ;
        RECT  0.140 0.520 1.180 0.680 ;
        RECT  0.940 0.520 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.250 1.760 5.390 1.920 ;
        RECT  1.020 0.520 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.230 1.760 5.390 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.250 1.760 4.410 2.100 ;
        RECT  2.780 1.940 4.410 2.100 ;
        RECT  5.950 1.200 6.110 2.100 ;
        RECT  5.230 1.940 6.110 2.100 ;
        RECT  3.340 0.300 4.410 0.460 ;
        RECT  5.230 0.300 6.750 0.460 ;
        RECT  4.250 0.300 4.410 0.640 ;
        RECT  5.230 0.300 5.390 0.640 ;
        RECT  4.250 0.480 5.390 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.590 0.300 6.750 1.160 ;
        RECT  6.590 1.000 7.130 1.160 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.070 0.640 6.430 0.800 ;
        RECT  12.010 1.120 12.530 1.280 ;
        RECT  8.750 1.520 9.590 1.680 ;
        RECT  10.070 1.520 10.910 1.680 ;
        RECT  12.010 1.120 12.170 1.740 ;
        RECT  11.390 1.580 12.170 1.740 ;
        RECT  7.430 1.700 8.270 1.860 ;
        RECT  6.270 0.640 6.430 2.100 ;
        RECT  8.110 1.700 8.270 2.100 ;
        RECT  9.430 1.520 9.590 2.100 ;
        RECT  10.750 1.520 10.910 2.100 ;
        RECT  7.430 1.700 7.590 2.100 ;
        RECT  6.270 1.940 7.590 2.100 ;
        RECT  8.750 1.520 8.910 2.100 ;
        RECT  8.110 1.940 8.910 2.100 ;
        RECT  10.070 1.520 10.230 2.100 ;
        RECT  9.430 1.940 10.230 2.100 ;
        RECT  11.390 1.580 11.550 2.100 ;
        RECT  10.750 1.940 11.550 2.100 ;
        RECT  12.590 0.620 12.870 0.960 ;
        RECT  11.510 0.800 12.870 0.960 ;
        RECT  11.510 0.800 11.670 1.360 ;
        RECT  12.690 0.620 12.870 1.900 ;
        RECT  12.390 1.700 12.870 1.900 ;
        RECT  9.260 0.300 10.230 0.460 ;
        RECT  10.750 0.300 11.670 0.460 ;
        RECT  12.270 0.300 13.190 0.460 ;
        RECT  11.510 0.300 11.670 0.640 ;
        RECT  10.070 0.300 10.230 0.700 ;
        RECT  12.270 0.300 12.430 0.640 ;
        RECT  11.510 0.480 12.430 0.640 ;
        RECT  7.020 0.480 8.590 0.680 ;
        RECT  10.750 0.300 10.910 0.700 ;
        RECT  10.070 0.540 10.910 0.700 ;
        RECT  13.030 0.300 13.190 1.260 ;
        RECT  9.260 0.300 9.420 1.200 ;
        RECT  8.430 1.040 9.420 1.200 ;
        RECT  13.030 1.100 14.670 1.260 ;
        RECT  7.070 1.380 8.590 1.540 ;
        RECT  7.070 1.380 7.270 1.780 ;
        RECT  8.430 0.480 8.590 1.780 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  4.130 1.140 5.090 2.400 ;
        RECT  0.000 1.160 5.090 2.400 ;
        RECT  6.700 1.140 16.000 2.400 ;
        RECT  0.000 1.200 16.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.000 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 16.000 1.140 ;
        RECT  3.400 0.000 4.130 1.160 ;
        RECT  5.090 0.000 6.700 1.200 ;
    END
END DFZRM8HM

MACRO DFZRM4HM
    CLASS CORE ;
    FOREIGN DFZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.620  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.430 0.620 8.700 1.200 ;
        RECT  8.430 0.620 8.590 1.760 ;
        RECT  8.310 0.620 8.700 0.840 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.210 1.440 11.900 1.640 ;
        RECT  11.700 0.720 11.900 1.640 ;
        RECT  11.210 0.720 11.900 0.920 ;
        RECT  11.210 1.440 11.410 2.080 ;
        RECT  11.210 0.440 11.410 0.920 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  11.730 1.840 11.930 2.540 ;
        RECT  10.600 1.480 10.800 2.540 ;
        RECT  9.070 1.840 9.270 2.540 ;
        RECT  7.750 2.020 7.950 2.540 ;
        RECT  4.790 2.080 5.070 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  11.730 -0.140 11.930 0.560 ;
        RECT  10.710 -0.140 10.870 0.760 ;
        RECT  9.190 -0.140 9.470 0.320 ;
        RECT  7.590 -0.140 7.790 0.560 ;
        RECT  4.790 -0.140 5.070 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.710 0.920 5.330 1.080 ;
        RECT  3.710 0.640 3.990 1.780 ;
        RECT  4.370 1.240 5.750 1.400 ;
        RECT  5.550 0.620 5.750 1.780 ;
        RECT  0.100 0.480 1.180 0.680 ;
        RECT  0.940 0.480 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.250 1.760 5.390 1.920 ;
        RECT  1.020 0.480 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.230 1.760 5.390 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.250 1.760 4.410 2.100 ;
        RECT  2.780 1.940 4.410 2.100 ;
        RECT  5.950 1.200 6.110 2.100 ;
        RECT  5.230 1.940 6.110 2.100 ;
        RECT  3.340 0.300 4.410 0.460 ;
        RECT  5.230 0.300 6.750 0.460 ;
        RECT  4.250 0.300 4.410 0.640 ;
        RECT  5.230 0.300 5.390 0.640 ;
        RECT  4.250 0.480 5.390 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.590 0.300 6.750 1.220 ;
        RECT  6.590 1.060 7.130 1.220 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.070 0.640 6.430 0.800 ;
        RECT  9.180 1.120 9.890 1.280 ;
        RECT  9.180 1.120 9.340 1.680 ;
        RECT  8.750 1.520 9.340 1.680 ;
        RECT  7.430 1.700 8.270 1.860 ;
        RECT  6.270 0.640 6.430 2.100 ;
        RECT  8.110 1.700 8.270 2.100 ;
        RECT  7.430 1.700 7.590 2.100 ;
        RECT  6.270 1.940 7.590 2.100 ;
        RECT  8.750 1.520 8.910 2.100 ;
        RECT  8.110 1.940 8.910 2.100 ;
        RECT  9.950 0.620 10.230 0.960 ;
        RECT  8.860 0.800 10.230 0.960 ;
        RECT  8.860 0.800 9.020 1.360 ;
        RECT  10.050 0.620 10.230 1.900 ;
        RECT  9.750 1.700 10.230 1.900 ;
        RECT  7.950 0.300 9.020 0.460 ;
        RECT  9.630 0.300 10.550 0.460 ;
        RECT  8.860 0.300 9.020 0.640 ;
        RECT  9.630 0.300 9.790 0.640 ;
        RECT  8.860 0.480 9.790 0.640 ;
        RECT  7.060 0.440 7.260 0.880 ;
        RECT  7.060 0.720 8.110 0.880 ;
        RECT  10.390 0.300 10.550 1.260 ;
        RECT  10.390 1.100 11.310 1.260 ;
        RECT  7.950 0.300 8.110 1.540 ;
        RECT  7.070 1.380 8.110 1.540 ;
        RECT  7.070 1.380 7.270 1.780 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  0.000 1.160 5.090 2.400 ;
        RECT  6.700 1.140 12.400 2.400 ;
        RECT  0.000 1.200 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 12.400 1.140 ;
        RECT  3.400 0.000 6.700 1.160 ;
        RECT  5.090 0.000 6.700 1.200 ;
    END
END DFZRM4HM

MACRO DFZRM2HM
    CLASS CORE ;
    FOREIGN DFZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.418  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.380 0.620 8.540 1.760 ;
        RECT  8.040 1.300 8.540 1.500 ;
        RECT  8.260 0.620 8.540 1.500 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.060 0.440 10.300 2.080 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.450 1.480 9.650 2.540 ;
        RECT  7.700 2.020 7.900 2.540 ;
        RECT  4.740 2.080 5.020 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.560 -0.140 9.720 0.760 ;
        RECT  7.500 -0.140 7.780 0.540 ;
        RECT  4.740 -0.140 5.020 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.660 0.920 5.280 1.080 ;
        RECT  3.660 0.640 3.940 1.780 ;
        RECT  4.320 1.240 5.700 1.400 ;
        RECT  5.500 0.620 5.700 1.780 ;
        RECT  0.100 0.480 1.180 0.680 ;
        RECT  0.940 0.480 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.200 1.760 5.340 1.920 ;
        RECT  1.020 0.480 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.180 1.760 5.340 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.200 1.760 4.360 2.100 ;
        RECT  2.780 1.940 4.360 2.100 ;
        RECT  5.900 1.200 6.060 2.100 ;
        RECT  5.180 1.940 6.060 2.100 ;
        RECT  3.340 0.300 4.360 0.460 ;
        RECT  5.180 0.300 6.700 0.460 ;
        RECT  4.200 0.300 4.360 0.640 ;
        RECT  5.180 0.300 5.340 0.640 ;
        RECT  4.200 0.480 5.340 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.540 0.300 6.700 1.220 ;
        RECT  6.540 1.060 7.080 1.220 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.020 0.640 6.380 0.800 ;
        RECT  7.380 1.700 8.220 1.860 ;
        RECT  6.220 0.640 6.380 2.100 ;
        RECT  8.060 1.700 8.220 2.100 ;
        RECT  7.380 1.700 7.540 2.100 ;
        RECT  6.220 1.940 7.540 2.100 ;
        RECT  8.060 1.940 8.780 2.100 ;
        RECT  8.720 1.040 9.080 1.320 ;
        RECT  8.800 0.620 9.080 1.660 ;
        RECT  7.940 0.300 9.400 0.460 ;
        RECT  7.010 0.320 7.210 0.880 ;
        RECT  7.940 0.300 8.100 0.880 ;
        RECT  7.010 0.720 8.100 0.880 ;
        RECT  9.240 0.300 9.400 1.260 ;
        RECT  9.240 1.100 9.780 1.260 ;
        RECT  7.300 0.720 7.460 1.540 ;
        RECT  7.020 1.380 7.460 1.540 ;
        RECT  7.020 1.380 7.220 1.780 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  0.000 1.160 5.040 2.400 ;
        RECT  6.650 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 10.400 1.140 ;
        RECT  3.400 0.000 6.650 1.160 ;
        RECT  5.040 0.000 6.650 1.200 ;
    END
END DFZRM2HM

MACRO DFZRM1HM
    CLASS CORE ;
    FOREIGN DFZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.314  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.380 0.620 8.540 1.760 ;
        RECT  8.040 1.300 8.540 1.500 ;
        RECT  8.260 0.620 8.540 1.500 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.060 0.520 10.300 1.810 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.450 1.530 9.650 2.540 ;
        RECT  7.700 2.020 7.900 2.540 ;
        RECT  4.740 2.080 5.020 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.560 -0.140 9.720 0.840 ;
        RECT  7.500 -0.140 7.780 0.540 ;
        RECT  4.740 -0.140 5.020 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.660 0.920 5.280 1.080 ;
        RECT  3.660 0.640 3.940 1.780 ;
        RECT  4.320 1.240 5.700 1.400 ;
        RECT  5.500 0.620 5.700 1.780 ;
        RECT  0.100 0.480 1.180 0.680 ;
        RECT  0.940 0.480 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.200 1.760 5.340 1.920 ;
        RECT  1.020 0.480 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.180 1.760 5.340 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.200 1.760 4.360 2.100 ;
        RECT  2.780 1.940 4.360 2.100 ;
        RECT  5.900 1.200 6.060 2.100 ;
        RECT  5.180 1.940 6.060 2.100 ;
        RECT  3.340 0.300 4.360 0.460 ;
        RECT  5.180 0.300 6.700 0.460 ;
        RECT  4.200 0.300 4.360 0.640 ;
        RECT  5.180 0.300 5.340 0.640 ;
        RECT  4.200 0.480 5.340 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.540 0.300 6.700 1.220 ;
        RECT  6.540 1.060 7.080 1.220 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.020 0.620 6.380 0.780 ;
        RECT  7.380 1.700 8.220 1.860 ;
        RECT  6.220 0.620 6.380 2.100 ;
        RECT  8.060 1.700 8.220 2.100 ;
        RECT  7.380 1.700 7.540 2.100 ;
        RECT  6.220 1.940 7.540 2.100 ;
        RECT  8.060 1.940 8.780 2.100 ;
        RECT  8.720 1.040 9.080 1.320 ;
        RECT  8.800 0.620 9.080 1.660 ;
        RECT  7.940 0.300 9.400 0.460 ;
        RECT  7.010 0.320 7.210 0.880 ;
        RECT  7.940 0.300 8.100 0.880 ;
        RECT  7.010 0.720 8.100 0.880 ;
        RECT  9.240 0.300 9.400 1.260 ;
        RECT  9.240 1.100 9.780 1.260 ;
        RECT  7.300 0.720 7.460 1.540 ;
        RECT  7.020 1.380 7.460 1.540 ;
        RECT  7.020 1.380 7.220 1.780 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  0.000 1.160 5.040 2.400 ;
        RECT  6.650 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 10.400 1.140 ;
        RECT  3.400 0.000 6.650 1.160 ;
        RECT  5.040 0.000 6.650 1.200 ;
    END
END DFZRM1HM

MACRO DFSM8HM
    CLASS CORE ;
    FOREIGN DFSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 13.562  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.080 7.100 1.280 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.770 1.020 7.460 1.340 ;
        RECT  7.300 0.300 7.460 1.340 ;
        RECT  5.350 0.300 7.460 0.460 ;
        RECT  4.800 1.020 5.520 1.300 ;
        RECT  5.350 0.300 5.520 1.300 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        ANTENNAGATEAREA 0.131  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.260  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.140 2.700 1.340 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.410 1.030 2.800 1.460 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.880 0.560 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.100 0.390 13.380 2.100 ;
        RECT  13.080 0.390 13.380 1.560 ;
        RECT  12.210 1.300 13.380 1.560 ;
        RECT  12.060 1.470 12.390 2.100 ;
        RECT  12.210 0.390 12.390 2.100 ;
        RECT  12.060 0.390 12.390 0.670 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.223  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.930 0.620 10.210 1.720 ;
        RECT  8.470 1.060 10.210 1.400 ;
        RECT  8.470 0.620 8.790 1.400 ;
        RECT  8.470 0.620 8.690 1.780 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.680 1.470 13.900 2.540 ;
        RECT  12.580 1.800 12.860 2.540 ;
        RECT  11.560 1.510 11.760 2.540 ;
        RECT  9.230 2.010 9.450 2.540 ;
        RECT  4.790 1.860 5.070 2.540 ;
        RECT  3.670 1.860 3.950 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.680 -0.140 13.900 0.670 ;
        RECT  12.580 -0.140 12.860 0.670 ;
        RECT  11.540 -0.140 11.820 0.780 ;
        RECT  9.290 -0.140 9.450 0.460 ;
        RECT  7.740 -0.140 7.960 0.580 ;
        RECT  3.670 -0.140 3.950 0.380 ;
        RECT  1.750 -0.140 2.050 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.400 0.920 0.680 ;
        RECT  0.740 0.990 1.640 1.240 ;
        RECT  0.740 0.400 0.920 1.920 ;
        RECT  0.100 1.720 0.920 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.290 2.100 ;
        RECT  2.730 0.640 3.120 0.840 ;
        RECT  2.960 0.640 3.120 1.780 ;
        RECT  2.960 0.900 4.170 1.060 ;
        RECT  3.880 0.900 4.170 1.260 ;
        RECT  2.960 0.900 3.150 1.780 ;
        RECT  2.500 1.620 3.150 1.780 ;
        RECT  2.330 0.300 3.510 0.460 ;
        RECT  4.150 0.300 5.190 0.460 ;
        RECT  4.910 0.300 5.190 0.500 ;
        RECT  3.350 0.300 3.510 0.720 ;
        RECT  4.150 0.300 4.310 0.720 ;
        RECT  3.350 0.550 4.310 0.720 ;
        RECT  1.150 0.530 2.510 0.760 ;
        RECT  2.330 0.300 2.510 0.790 ;
        RECT  1.870 0.530 2.510 0.790 ;
        RECT  1.870 0.530 2.150 1.600 ;
        RECT  1.110 1.400 2.150 1.600 ;
        RECT  4.470 0.640 4.830 0.840 ;
        RECT  3.370 1.240 3.670 1.700 ;
        RECT  4.470 0.640 4.640 1.700 ;
        RECT  3.370 1.540 5.550 1.700 ;
        RECT  5.270 1.540 5.550 1.850 ;
        RECT  6.260 0.620 7.140 0.840 ;
        RECT  8.000 1.060 8.300 1.340 ;
        RECT  6.260 0.620 6.420 1.780 ;
        RECT  8.000 1.060 8.210 1.780 ;
        RECT  6.260 1.580 8.210 1.780 ;
        RECT  5.690 0.640 6.060 0.920 ;
        RECT  10.370 1.090 10.960 1.310 ;
        RECT  8.910 1.610 9.770 1.770 ;
        RECT  9.610 1.610 9.770 2.040 ;
        RECT  5.900 0.640 6.060 2.100 ;
        RECT  10.370 1.090 10.530 2.040 ;
        RECT  9.610 1.880 10.530 2.040 ;
        RECT  8.910 1.610 9.070 2.100 ;
        RECT  5.900 1.940 9.070 2.100 ;
        RECT  8.130 0.300 9.110 0.460 ;
        RECT  9.610 0.300 10.530 0.460 ;
        RECT  8.950 0.300 9.110 0.810 ;
        RECT  10.370 0.300 10.530 0.920 ;
        RECT  9.610 0.300 9.770 0.810 ;
        RECT  8.950 0.650 9.770 0.810 ;
        RECT  8.130 0.300 8.290 0.900 ;
        RECT  7.620 0.740 8.290 0.900 ;
        RECT  11.020 0.500 11.300 0.920 ;
        RECT  10.370 0.760 11.300 0.920 ;
        RECT  7.620 0.740 7.840 1.240 ;
        RECT  11.130 0.960 12.000 1.300 ;
        RECT  11.130 0.500 11.300 1.740 ;
        RECT  11.080 1.440 11.300 1.740 ;
        LAYER VTPH ;
        RECT  0.530 1.080 1.990 2.400 ;
        RECT  0.000 1.140 2.150 2.400 ;
        RECT  3.570 1.160 5.310 2.400 ;
        RECT  0.000 1.200 5.310 2.400 ;
        RECT  6.750 1.140 14.000 2.400 ;
        RECT  0.000 1.240 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 0.530 1.140 ;
        RECT  1.990 0.000 14.000 1.140 ;
        RECT  2.150 0.000 6.750 1.160 ;
        RECT  2.150 0.000 3.570 1.200 ;
        RECT  5.310 0.000 6.750 1.240 ;
    END
END DFSM8HM

MACRO DFSM4HM
    CLASS CORE ;
    FOREIGN DFSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        ANTENNAGATEAREA 0.124  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.450  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.420 1.140 2.620 1.340 ;
        LAYER ME2 ;
        RECT  2.420 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.330 1.030 2.720 1.460 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 13.562  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.080 7.100 1.280 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.690 1.020 7.380 1.340 ;
        RECT  7.220 0.300 7.380 1.340 ;
        RECT  5.270 0.300 7.380 0.460 ;
        RECT  4.720 1.020 5.440 1.300 ;
        RECT  5.270 0.300 5.440 1.300 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.380 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.430 0.840 11.160 1.560 ;
        RECT  10.430 0.390 10.710 2.100 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.392  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.390 0.620 8.760 1.780 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.950 1.800 11.230 2.540 ;
        RECT  9.910 1.600 10.190 2.540 ;
        RECT  4.710 1.860 4.990 2.540 ;
        RECT  3.590 1.860 3.870 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.950 -0.140 11.230 0.670 ;
        RECT  9.910 -0.140 10.190 0.780 ;
        RECT  7.660 -0.140 7.880 0.580 ;
        RECT  3.590 -0.140 3.870 0.380 ;
        RECT  1.670 -0.140 1.970 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.920 0.560 ;
        RECT  0.740 0.990 1.260 1.240 ;
        RECT  0.740 0.300 0.920 1.920 ;
        RECT  0.100 1.590 0.920 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.210 2.100 ;
        RECT  2.650 0.640 3.040 0.840 ;
        RECT  2.880 0.640 3.040 1.780 ;
        RECT  2.880 0.900 4.090 1.060 ;
        RECT  3.800 0.900 4.090 1.260 ;
        RECT  2.880 0.900 3.070 1.780 ;
        RECT  2.420 1.620 3.070 1.780 ;
        RECT  2.250 0.300 3.430 0.460 ;
        RECT  4.070 0.300 5.110 0.460 ;
        RECT  4.830 0.300 5.110 0.500 ;
        RECT  3.270 0.300 3.430 0.720 ;
        RECT  4.070 0.300 4.230 0.720 ;
        RECT  3.270 0.550 4.230 0.720 ;
        RECT  2.250 0.300 2.430 0.760 ;
        RECT  1.150 0.530 2.430 0.760 ;
        RECT  1.790 0.530 2.070 1.600 ;
        RECT  1.110 1.400 2.070 1.600 ;
        RECT  4.390 0.640 4.750 0.840 ;
        RECT  3.290 1.240 3.590 1.700 ;
        RECT  4.390 0.640 4.560 1.700 ;
        RECT  3.290 1.540 5.470 1.700 ;
        RECT  5.190 1.540 5.470 1.850 ;
        RECT  6.180 0.620 7.060 0.840 ;
        RECT  6.180 0.620 6.340 1.780 ;
        RECT  7.960 1.060 8.220 1.780 ;
        RECT  6.180 1.580 8.220 1.780 ;
        RECT  5.610 0.640 5.980 0.920 ;
        RECT  5.820 0.640 5.980 2.100 ;
        RECT  9.130 1.010 9.290 2.100 ;
        RECT  5.820 1.940 9.290 2.100 ;
        RECT  8.050 0.300 9.670 0.460 ;
        RECT  8.050 0.300 8.210 0.900 ;
        RECT  7.540 0.740 8.210 0.900 ;
        RECT  7.540 0.740 7.760 1.240 ;
        RECT  9.450 0.960 10.270 1.240 ;
        RECT  9.450 0.300 9.670 1.740 ;
        LAYER VTPH ;
        RECT  0.530 1.080 1.910 2.400 ;
        RECT  0.000 1.140 2.070 2.400 ;
        RECT  3.490 1.160 5.230 2.400 ;
        RECT  0.000 1.200 5.230 2.400 ;
        RECT  6.670 1.140 11.600 2.400 ;
        RECT  0.000 1.240 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.080 ;
        RECT  0.000 0.000 0.530 1.140 ;
        RECT  1.910 0.000 11.600 1.140 ;
        RECT  2.070 0.000 6.670 1.160 ;
        RECT  2.070 0.000 3.490 1.200 ;
        RECT  5.230 0.000 6.670 1.240 ;
    END
END DFSM4HM

MACRO DFSM2HM
    CLASS CORE ;
    FOREIGN DFSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.356  LAYER ME1  ;
        ANTENNADIFFAREA 0.356  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.450 0.660 8.650 0.860 ;
        LAYER ME2 ;
        RECT  8.450 0.420 8.700 1.160 ;
        LAYER ME1 ;
        RECT  8.350 0.620 8.720 0.920 ;
        RECT  8.290 1.440 8.510 1.740 ;
        RECT  8.350 0.620 8.510 1.740 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        ANTENNAGATEAREA 0.124  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.450  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.390 1.140 2.590 1.340 ;
        LAYER ME2 ;
        RECT  2.390 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.290 1.030 2.680 1.460 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.450 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.080 0.300 10.300 2.100 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        ANTENNAGATEAREA 0.196  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 13.532  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.080 7.100 1.280 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.670 1.020 7.360 1.340 ;
        RECT  7.200 0.300 7.360 1.340 ;
        RECT  5.230 0.300 7.360 0.460 ;
        RECT  4.680 1.020 5.390 1.300 ;
        RECT  5.230 0.300 5.390 1.300 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.500 1.820 9.780 2.540 ;
        RECT  4.670 1.860 4.950 2.540 ;
        RECT  3.550 1.860 3.830 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.500 -0.140 9.780 0.500 ;
        RECT  7.640 -0.140 7.860 0.580 ;
        RECT  3.550 -0.140 3.830 0.380 ;
        RECT  1.620 -0.140 1.920 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.400 0.830 0.680 ;
        RECT  0.650 0.920 1.200 1.120 ;
        RECT  0.650 0.400 0.830 1.920 ;
        RECT  0.100 1.720 0.830 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.170 2.100 ;
        RECT  2.610 0.640 3.020 0.840 ;
        RECT  2.840 0.640 3.020 1.780 ;
        RECT  2.840 0.900 4.050 1.060 ;
        RECT  3.760 0.900 4.050 1.200 ;
        RECT  2.840 0.900 3.030 1.780 ;
        RECT  2.410 1.620 3.030 1.780 ;
        RECT  2.210 0.300 3.390 0.460 ;
        RECT  4.030 0.300 5.070 0.460 ;
        RECT  4.790 0.300 5.070 0.500 ;
        RECT  3.230 0.300 3.390 0.720 ;
        RECT  2.210 0.300 2.390 0.720 ;
        RECT  1.020 0.530 2.390 0.720 ;
        RECT  4.030 0.300 4.190 0.720 ;
        RECT  3.230 0.550 4.190 0.720 ;
        RECT  1.020 0.530 2.030 0.740 ;
        RECT  1.870 0.530 2.030 1.600 ;
        RECT  1.050 1.400 2.030 1.600 ;
        RECT  4.350 0.640 4.710 0.840 ;
        RECT  3.250 1.240 3.470 1.700 ;
        RECT  4.350 0.640 4.520 1.700 ;
        RECT  3.250 1.540 5.430 1.700 ;
        RECT  5.150 1.540 5.430 1.810 ;
        RECT  6.160 0.620 7.040 0.840 ;
        RECT  7.940 1.060 8.160 1.340 ;
        RECT  6.160 0.620 6.320 1.740 ;
        RECT  7.940 1.060 8.100 1.740 ;
        RECT  6.160 1.580 8.100 1.740 ;
        RECT  5.560 0.640 5.900 0.860 ;
        RECT  8.670 1.120 9.320 1.280 ;
        RECT  5.740 0.640 5.900 2.060 ;
        RECT  8.670 1.120 8.830 2.060 ;
        RECT  5.740 1.900 8.830 2.060 ;
        RECT  8.030 0.300 9.220 0.460 ;
        RECT  9.000 0.300 9.220 0.840 ;
        RECT  9.000 0.660 9.920 0.840 ;
        RECT  8.030 0.300 8.190 0.900 ;
        RECT  7.520 0.740 8.190 0.900 ;
        RECT  7.520 0.740 7.740 1.240 ;
        RECT  9.700 0.660 9.920 1.660 ;
        RECT  9.000 1.500 9.920 1.660 ;
        RECT  9.000 1.500 9.220 1.830 ;
        LAYER VTPH ;
        RECT  0.530 1.080 1.950 2.400 ;
        RECT  0.000 1.140 1.950 2.400 ;
        RECT  3.450 1.160 5.100 2.400 ;
        RECT  6.630 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 0.530 1.140 ;
        RECT  1.950 0.000 10.400 1.140 ;
        RECT  1.950 0.000 6.630 1.160 ;
        RECT  1.950 0.000 3.450 1.200 ;
        RECT  5.100 0.000 6.630 1.200 ;
    END
END DFSM2HM

MACRO DFSM1HM
    CLASS CORE ;
    FOREIGN DFSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.281  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.390 1.140 2.590 1.340 ;
        LAYER ME2 ;
        RECT  2.390 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.290 1.030 2.680 1.460 ;
        END
    END D
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.291  LAYER ME1  ;
        ANTENNADIFFAREA 0.291  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.450 0.660 8.650 0.860 ;
        LAYER ME2 ;
        RECT  8.450 0.420 8.700 1.160 ;
        LAYER ME1 ;
        RECT  8.350 0.620 8.720 0.920 ;
        RECT  8.290 1.440 8.510 1.740 ;
        RECT  8.350 0.620 8.510 1.740 ;
        END
    END QB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.068  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 0.450 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.282  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.080 0.300 10.300 2.050 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        ANTENNAGATEAREA 0.152  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 17.367  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.080 7.100 1.280 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.670 1.020 7.360 1.340 ;
        RECT  7.200 0.300 7.360 1.340 ;
        RECT  5.230 0.300 7.360 0.460 ;
        RECT  4.680 1.020 5.390 1.300 ;
        RECT  5.230 0.300 5.390 1.300 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.500 1.760 9.780 2.540 ;
        RECT  4.670 1.860 4.950 2.540 ;
        RECT  3.550 1.860 3.830 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.500 -0.140 9.780 0.500 ;
        RECT  7.640 -0.140 7.860 0.560 ;
        RECT  3.550 -0.140 3.830 0.380 ;
        RECT  1.620 -0.140 1.920 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.400 0.830 0.680 ;
        RECT  0.650 0.920 1.200 1.120 ;
        RECT  0.650 0.400 0.830 1.920 ;
        RECT  0.100 1.720 0.830 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.170 2.100 ;
        RECT  2.610 0.640 3.020 0.840 ;
        RECT  2.840 0.640 3.020 1.780 ;
        RECT  2.840 0.900 4.050 1.060 ;
        RECT  3.760 0.900 4.050 1.200 ;
        RECT  2.840 0.900 3.030 1.780 ;
        RECT  2.410 1.620 3.030 1.780 ;
        RECT  2.210 0.300 3.390 0.460 ;
        RECT  4.030 0.300 5.070 0.460 ;
        RECT  4.790 0.300 5.070 0.500 ;
        RECT  3.230 0.300 3.390 0.720 ;
        RECT  2.210 0.300 2.390 0.720 ;
        RECT  1.020 0.530 2.390 0.720 ;
        RECT  4.030 0.300 4.190 0.720 ;
        RECT  3.230 0.550 4.190 0.720 ;
        RECT  1.020 0.530 2.030 0.740 ;
        RECT  1.870 0.530 2.030 1.600 ;
        RECT  1.050 1.400 2.030 1.600 ;
        RECT  4.350 0.640 4.710 0.840 ;
        RECT  3.250 1.240 3.470 1.700 ;
        RECT  4.350 0.640 4.520 1.700 ;
        RECT  3.250 1.540 5.430 1.700 ;
        RECT  5.150 1.540 5.430 1.810 ;
        RECT  6.160 0.620 7.040 0.840 ;
        RECT  7.940 1.060 8.160 1.340 ;
        RECT  6.160 0.620 6.320 1.740 ;
        RECT  7.940 1.060 8.100 1.740 ;
        RECT  6.160 1.580 8.100 1.740 ;
        RECT  5.560 0.640 5.900 0.860 ;
        RECT  8.670 1.120 9.320 1.280 ;
        RECT  5.740 0.640 5.900 2.060 ;
        RECT  8.670 1.120 8.830 2.060 ;
        RECT  5.740 1.900 8.830 2.060 ;
        RECT  8.030 0.300 9.220 0.460 ;
        RECT  9.000 0.300 9.220 0.840 ;
        RECT  9.000 0.660 9.920 0.840 ;
        RECT  8.030 0.300 8.190 0.900 ;
        RECT  7.520 0.740 8.190 0.900 ;
        RECT  7.520 0.740 7.740 1.240 ;
        RECT  9.700 0.660 9.920 1.600 ;
        RECT  9.000 1.440 9.920 1.600 ;
        RECT  9.000 1.440 9.220 1.830 ;
        LAYER VTPH ;
        RECT  0.530 1.080 1.950 2.400 ;
        RECT  0.000 1.140 1.950 2.400 ;
        RECT  3.450 1.160 5.100 2.400 ;
        RECT  6.630 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 0.530 1.140 ;
        RECT  1.950 0.000 10.400 1.140 ;
        RECT  1.950 0.000 6.630 1.160 ;
        RECT  1.950 0.000 3.450 1.200 ;
        RECT  5.100 0.000 6.630 1.200 ;
    END
END DFSM1HM

MACRO DFRSM8HM
    CLASS CORE ;
    FOREIGN DFRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.112  LAYER ME1  ;
        ANTENNAGATEAREA 0.112  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 17.892  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.160 1.650 9.360 1.850 ;
        LAYER ME2 ;
        RECT  9.160 1.240 9.500 1.960 ;
        LAYER ME1 ;
        RECT  6.360 1.920 9.360 2.080 ;
        RECT  9.160 1.500 9.360 2.080 ;
        RECT  6.360 1.660 6.520 2.080 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.570 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.380 1.380 14.860 1.600 ;
        RECT  13.420 0.680 14.820 0.840 ;
        RECT  14.520 0.380 14.820 0.840 ;
        RECT  14.040 0.680 14.360 1.600 ;
        RECT  13.420 0.380 13.700 0.840 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.981  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.700 0.380 16.980 2.100 ;
        RECT  15.660 0.840 16.980 1.160 ;
        RECT  15.660 0.380 15.940 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.259  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.080 0.900 12.820 1.180 ;
        RECT  12.080 0.300 12.260 1.180 ;
        RECT  10.510 0.300 12.260 0.460 ;
        RECT  10.270 0.500 10.680 0.870 ;
        RECT  10.510 0.300 10.680 0.870 ;
        RECT  9.350 0.500 10.680 0.710 ;
        RECT  9.350 0.300 9.510 0.710 ;
        RECT  8.180 0.300 9.510 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.600 2.540 ;
        RECT  17.220 1.500 17.500 2.540 ;
        RECT  16.180 1.480 16.450 2.540 ;
        RECT  15.100 2.080 15.380 2.540 ;
        RECT  13.980 2.080 14.260 2.540 ;
        RECT  12.860 2.080 13.140 2.540 ;
        RECT  10.560 1.760 10.780 2.540 ;
        RECT  9.520 1.860 9.800 2.540 ;
        RECT  5.980 1.730 6.140 2.540 ;
        RECT  4.720 1.800 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.600 0.140 ;
        RECT  17.220 -0.140 17.500 0.660 ;
        RECT  16.180 -0.140 16.450 0.660 ;
        RECT  15.100 -0.140 15.380 0.660 ;
        RECT  13.980 -0.140 14.260 0.520 ;
        RECT  12.820 -0.140 13.100 0.660 ;
        RECT  10.020 -0.140 10.300 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.400 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.720 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.640 ;
        RECT  4.200 1.440 5.260 1.640 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  4.520 1.120 5.620 1.280 ;
        RECT  6.240 0.620 6.520 1.500 ;
        RECT  5.420 1.340 6.960 1.500 ;
        RECT  6.680 1.340 6.960 1.760 ;
        RECT  5.420 1.120 5.620 1.800 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 7.000 0.460 ;
        RECT  1.150 0.330 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.790 0.300 7.000 1.180 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.070 1.440 2.070 1.600 ;
        RECT  7.260 0.520 7.420 1.760 ;
        RECT  7.260 0.880 8.680 1.160 ;
        RECT  7.260 0.880 7.520 1.760 ;
        RECT  7.160 1.600 7.520 1.760 ;
        RECT  13.010 1.000 13.620 1.160 ;
        RECT  9.860 1.060 11.920 1.260 ;
        RECT  11.640 0.620 11.920 1.600 ;
        RECT  11.260 1.060 11.920 1.600 ;
        RECT  13.010 1.000 13.170 1.600 ;
        RECT  11.260 1.370 13.170 1.600 ;
        RECT  11.260 1.060 11.580 1.660 ;
        RECT  8.840 0.620 9.150 1.250 ;
        RECT  15.040 0.960 15.480 1.240 ;
        RECT  8.840 1.090 9.700 1.250 ;
        RECT  9.540 1.090 9.700 1.660 ;
        RECT  9.540 1.420 11.100 1.580 ;
        RECT  9.540 1.420 10.400 1.660 ;
        RECT  8.840 0.620 9.000 1.740 ;
        RECT  7.800 1.540 9.000 1.740 ;
        RECT  10.940 1.420 11.100 1.980 ;
        RECT  11.710 1.760 15.240 1.920 ;
        RECT  15.040 0.960 15.240 1.920 ;
        RECT  10.940 1.820 11.870 1.980 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.630 2.400 ;
        RECT  10.380 1.080 11.450 2.400 ;
        RECT  12.100 1.080 15.470 2.400 ;
        RECT  0.000 1.140 7.090 2.400 ;
        RECT  8.080 1.140 17.600 2.400 ;
        RECT  0.000 1.200 17.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.600 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.630 0.000 10.380 1.140 ;
        RECT  11.450 0.000 12.100 1.140 ;
        RECT  15.550 0.000 17.600 1.140 ;
        RECT  7.090 0.000 8.080 1.200 ;
    END
END DFRSM8HM

MACRO DFRSM4HM
    CLASS CORE ;
    FOREIGN DFRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.112  LAYER ME1  ;
        ANTENNAGATEAREA 0.112  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 17.892  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.160 1.650 9.360 1.850 ;
        LAYER ME2 ;
        RECT  9.160 1.240 9.500 1.960 ;
        LAYER ME1 ;
        RECT  6.360 1.920 9.360 2.080 ;
        RECT  9.160 1.500 9.360 2.080 ;
        RECT  6.360 1.660 6.520 2.080 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.570 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.380 1.380 13.910 1.600 ;
        RECT  13.590 0.680 13.910 1.600 ;
        RECT  13.420 0.380 13.700 0.840 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.485  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.540 0.840 15.100 1.160 ;
        RECT  14.540 0.380 14.820 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.260  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.080 0.900 12.820 1.180 ;
        RECT  12.080 0.300 12.260 1.180 ;
        RECT  10.510 0.300 12.260 0.460 ;
        RECT  10.270 0.500 10.680 0.870 ;
        RECT  10.510 0.300 10.680 0.870 ;
        RECT  9.350 0.500 10.680 0.710 ;
        RECT  9.350 0.300 9.510 0.710 ;
        RECT  8.180 0.300 9.510 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  15.060 1.480 15.340 2.540 ;
        RECT  13.980 2.080 14.260 2.540 ;
        RECT  12.860 2.080 13.140 2.540 ;
        RECT  10.560 1.760 10.780 2.540 ;
        RECT  9.520 1.860 9.800 2.540 ;
        RECT  5.980 1.730 6.140 2.540 ;
        RECT  4.720 1.800 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  15.060 -0.140 15.340 0.660 ;
        RECT  13.980 -0.140 14.260 0.520 ;
        RECT  12.820 -0.140 13.100 0.660 ;
        RECT  10.020 -0.140 10.300 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.260 1.260 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.720 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.640 ;
        RECT  4.200 1.440 5.260 1.640 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  4.520 1.120 5.620 1.280 ;
        RECT  6.240 0.620 6.520 1.500 ;
        RECT  5.420 1.340 6.960 1.500 ;
        RECT  6.680 1.340 6.960 1.760 ;
        RECT  5.420 1.120 5.620 1.800 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 7.000 0.460 ;
        RECT  1.150 0.330 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.790 0.300 7.000 1.180 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.070 1.440 2.070 1.600 ;
        RECT  7.220 0.520 7.380 1.760 ;
        RECT  7.220 0.880 8.680 1.160 ;
        RECT  7.220 0.880 7.520 1.760 ;
        RECT  7.160 1.600 7.520 1.760 ;
        RECT  13.010 1.000 13.430 1.160 ;
        RECT  9.860 1.060 11.920 1.260 ;
        RECT  11.640 0.620 11.920 1.600 ;
        RECT  11.260 1.060 11.920 1.600 ;
        RECT  13.010 1.000 13.170 1.600 ;
        RECT  11.260 1.370 13.170 1.600 ;
        RECT  11.260 1.060 11.580 1.660 ;
        RECT  8.840 0.620 9.150 1.250 ;
        RECT  14.120 0.960 14.360 1.240 ;
        RECT  8.840 1.090 9.700 1.250 ;
        RECT  9.540 1.090 9.700 1.660 ;
        RECT  9.540 1.420 11.100 1.580 ;
        RECT  9.540 1.420 10.400 1.660 ;
        RECT  8.840 0.620 9.000 1.740 ;
        RECT  7.800 1.540 9.000 1.740 ;
        RECT  10.940 1.420 11.100 1.980 ;
        RECT  11.710 1.760 14.320 1.920 ;
        RECT  14.120 0.960 14.320 1.920 ;
        RECT  10.940 1.820 11.870 1.980 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.630 2.400 ;
        RECT  10.380 1.080 11.450 2.400 ;
        RECT  12.100 1.080 14.430 2.400 ;
        RECT  0.000 1.140 7.050 2.400 ;
        RECT  8.080 1.140 15.600 2.400 ;
        RECT  0.000 1.200 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.630 0.000 10.380 1.140 ;
        RECT  11.450 0.000 12.100 1.140 ;
        RECT  14.430 0.000 15.600 1.140 ;
        RECT  7.050 0.000 8.080 1.200 ;
    END
END DFRSM4HM

MACRO DFRSM2HM
    CLASS CORE ;
    FOREIGN DFRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        ANTENNAGATEAREA 0.096  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 20.800  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.160 1.650 9.360 1.850 ;
        LAYER ME2 ;
        RECT  9.160 1.240 9.500 1.960 ;
        LAYER ME1 ;
        RECT  6.360 1.920 9.360 2.080 ;
        RECT  9.160 1.500 9.360 2.080 ;
        RECT  6.360 1.660 6.520 2.080 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.440 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.430 1.400 12.790 1.600 ;
        RECT  12.500 0.380 12.790 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.570 0.380 13.900 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.330 0.500 10.690 0.870 ;
        RECT  9.350 0.500 10.690 0.710 ;
        RECT  9.350 0.300 9.510 0.710 ;
        RECT  8.180 0.300 9.510 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  12.950 2.080 13.230 2.540 ;
        RECT  11.840 2.080 12.120 2.540 ;
        RECT  10.580 1.800 10.800 2.540 ;
        RECT  9.520 1.860 9.800 2.540 ;
        RECT  5.980 1.730 6.140 2.540 ;
        RECT  4.720 1.800 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  12.970 -0.140 13.250 0.520 ;
        RECT  12.010 -0.140 12.170 0.700 ;
        RECT  10.020 -0.140 10.300 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.720 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.640 ;
        RECT  4.200 1.440 5.260 1.640 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  4.520 1.120 5.620 1.280 ;
        RECT  6.240 0.620 6.520 1.500 ;
        RECT  5.420 1.340 6.960 1.500 ;
        RECT  6.680 1.340 6.960 1.760 ;
        RECT  5.420 1.120 5.620 1.800 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 7.000 0.460 ;
        RECT  1.150 0.350 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.790 0.300 7.000 1.180 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.100 1.440 2.070 1.600 ;
        RECT  7.260 0.520 7.420 1.760 ;
        RECT  7.260 0.880 8.680 1.160 ;
        RECT  7.260 0.880 7.520 1.760 ;
        RECT  7.160 1.600 7.520 1.760 ;
        RECT  11.460 0.500 11.740 1.220 ;
        RECT  11.460 1.000 12.330 1.220 ;
        RECT  9.860 1.060 11.560 1.260 ;
        RECT  11.280 1.060 11.560 1.600 ;
        RECT  8.840 0.620 9.150 1.250 ;
        RECT  8.840 1.090 9.700 1.250 ;
        RECT  9.540 1.090 9.700 1.660 ;
        RECT  9.540 1.420 11.120 1.580 ;
        RECT  9.540 1.420 10.360 1.660 ;
        RECT  8.840 0.620 9.000 1.740 ;
        RECT  7.800 1.540 9.000 1.740 ;
        RECT  10.960 1.420 11.120 1.920 ;
        RECT  13.160 0.960 13.390 1.920 ;
        RECT  10.960 1.760 13.390 1.920 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.630 2.400 ;
        RECT  10.380 1.080 12.940 2.400 ;
        RECT  0.000 1.140 7.090 2.400 ;
        RECT  8.080 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.630 0.000 10.380 1.140 ;
        RECT  12.940 0.000 14.000 1.140 ;
        RECT  7.090 0.000 8.080 1.200 ;
    END
END DFRSM2HM

MACRO DFRSM1HM
    CLASS CORE ;
    FOREIGN DFRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.655  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 23.111  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  9.160 1.650 9.360 1.850 ;
        LAYER ME2 ;
        RECT  9.160 1.240 9.500 1.960 ;
        LAYER ME1 ;
        RECT  6.360 1.920 9.360 2.080 ;
        RECT  9.160 1.500 9.360 2.080 ;
        RECT  6.360 1.660 6.520 2.080 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.440 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.430 1.400 12.790 1.600 ;
        RECT  12.500 0.380 12.790 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.570 0.380 13.900 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.330 0.500 10.690 0.870 ;
        RECT  9.350 0.500 10.690 0.710 ;
        RECT  9.350 0.300 9.510 0.710 ;
        RECT  8.180 0.300 9.510 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  12.950 2.080 13.230 2.540 ;
        RECT  11.840 2.080 12.120 2.540 ;
        RECT  10.580 1.800 10.800 2.540 ;
        RECT  9.520 1.860 9.800 2.540 ;
        RECT  5.980 1.730 6.140 2.540 ;
        RECT  4.720 1.800 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  12.970 -0.140 13.250 0.520 ;
        RECT  12.010 -0.140 12.170 0.700 ;
        RECT  10.020 -0.140 10.300 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.720 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.640 ;
        RECT  4.200 1.440 5.260 1.640 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  4.520 1.120 5.620 1.280 ;
        RECT  6.240 0.620 6.520 1.500 ;
        RECT  5.420 1.340 6.960 1.500 ;
        RECT  6.680 1.340 6.960 1.760 ;
        RECT  5.420 1.120 5.620 1.790 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 7.000 0.460 ;
        RECT  1.150 0.350 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.790 0.300 7.000 1.180 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.100 1.440 2.070 1.600 ;
        RECT  7.260 0.520 7.420 1.760 ;
        RECT  7.260 0.880 8.680 1.160 ;
        RECT  7.260 0.880 7.520 1.760 ;
        RECT  7.160 1.600 7.520 1.760 ;
        RECT  11.460 0.340 11.740 1.220 ;
        RECT  11.460 1.000 12.330 1.220 ;
        RECT  9.860 1.060 11.560 1.260 ;
        RECT  11.280 1.060 11.560 1.600 ;
        RECT  8.840 0.620 9.150 1.250 ;
        RECT  8.840 1.090 9.700 1.250 ;
        RECT  9.540 1.090 9.700 1.660 ;
        RECT  9.540 1.420 11.120 1.580 ;
        RECT  9.540 1.420 10.360 1.660 ;
        RECT  8.840 0.620 9.000 1.740 ;
        RECT  7.800 1.540 9.000 1.740 ;
        RECT  10.960 1.420 11.120 1.920 ;
        RECT  13.160 0.960 13.390 1.920 ;
        RECT  10.960 1.760 13.390 1.920 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.630 2.400 ;
        RECT  10.380 1.080 12.940 2.400 ;
        RECT  0.000 1.140 7.090 2.400 ;
        RECT  8.080 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.630 0.000 10.380 1.140 ;
        RECT  12.940 0.000 14.000 1.140 ;
        RECT  7.090 0.000 8.080 1.200 ;
    END
END DFRSM1HM

MACRO DFRM8HM
    CLASS CORE ;
    FOREIGN DFRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.570 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.670 1.330 13.160 1.600 ;
        RECT  12.860 0.380 13.160 1.600 ;
        RECT  11.640 0.680 13.160 0.840 ;
        RECT  12.810 0.380 13.160 0.840 ;
        RECT  11.640 0.300 11.960 0.840 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.981  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.980 0.380 15.270 2.100 ;
        RECT  13.950 1.220 15.270 1.560 ;
        RECT  13.950 0.380 14.250 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.510 0.900 11.110 1.180 ;
        RECT  10.510 0.300 10.710 1.180 ;
        RECT  9.220 0.300 10.710 0.460 ;
        RECT  8.160 0.500 9.390 0.870 ;
        RECT  9.220 0.300 9.390 0.870 ;
        RECT  8.160 0.300 8.320 0.870 ;
        RECT  7.300 0.300 8.320 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.000 2.540 ;
        RECT  15.510 1.500 15.790 2.540 ;
        RECT  14.470 1.840 14.740 2.540 ;
        RECT  13.390 2.080 13.670 2.540 ;
        RECT  12.270 2.080 12.550 2.540 ;
        RECT  10.020 2.080 10.300 2.540 ;
        RECT  8.600 1.860 8.880 2.540 ;
        RECT  4.780 1.760 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.000 0.140 ;
        RECT  15.510 -0.140 15.790 0.660 ;
        RECT  14.470 -0.140 14.740 0.660 ;
        RECT  13.390 -0.140 13.670 0.660 ;
        RECT  12.270 -0.140 12.550 0.520 ;
        RECT  11.110 -0.140 11.390 0.660 ;
        RECT  8.640 -0.140 8.920 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.400 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.720 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.600 ;
        RECT  4.200 1.440 5.330 1.600 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  5.170 1.440 5.330 2.020 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  5.860 0.620 6.200 1.280 ;
        RECT  4.520 1.120 6.200 1.280 ;
        RECT  5.490 1.120 5.710 1.960 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 6.540 0.460 ;
        RECT  1.150 0.330 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.380 0.300 6.540 1.330 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.070 1.440 2.070 1.600 ;
        RECT  6.700 0.950 7.560 1.230 ;
        RECT  6.700 0.560 6.860 1.960 ;
        RECT  6.070 1.640 6.860 1.960 ;
        RECT  11.300 1.000 12.670 1.160 ;
        RECT  8.160 1.100 10.350 1.320 ;
        RECT  10.070 0.620 10.350 1.600 ;
        RECT  9.360 1.100 10.350 1.600 ;
        RECT  11.300 1.000 11.460 1.600 ;
        RECT  9.360 1.370 11.460 1.600 ;
        RECT  13.330 0.960 13.770 1.240 ;
        RECT  7.720 0.620 8.000 1.960 ;
        RECT  7.020 1.520 8.000 1.960 ;
        RECT  7.020 1.540 9.200 1.700 ;
        RECT  9.040 1.540 9.200 1.920 ;
        RECT  13.330 0.960 13.530 1.920 ;
        RECT  9.040 1.760 13.530 1.920 ;
        RECT  7.020 1.540 8.200 1.960 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.630 2.400 ;
        RECT  9.120 1.080 9.880 2.400 ;
        RECT  10.530 1.080 13.840 2.400 ;
        RECT  0.000 1.140 5.900 2.400 ;
        RECT  7.910 1.140 16.000 2.400 ;
        RECT  0.000 1.260 16.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.000 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.630 0.000 9.120 1.140 ;
        RECT  9.880 0.000 10.530 1.140 ;
        RECT  13.840 0.000 16.000 1.140 ;
        RECT  5.900 0.000 7.910 1.260 ;
    END
END DFRM8HM

MACRO DFRM4HM
    CLASS CORE ;
    FOREIGN DFRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.318  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.200 1.100 0.400 1.300 ;
        LAYER ME2 ;
        RECT  0.100 0.900 0.430 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.020 0.570 1.360 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.670 1.330 12.300 1.600 ;
        RECT  12.090 0.680 12.300 1.600 ;
        RECT  11.640 0.680 12.300 0.840 ;
        RECT  11.640 0.300 11.960 0.840 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.485  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.890 1.480 13.630 1.680 ;
        RECT  13.470 0.720 13.630 1.680 ;
        RECT  12.830 0.720 13.630 0.880 ;
        RECT  12.890 1.480 13.180 2.100 ;
        RECT  12.830 0.380 13.180 0.880 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.510 0.900 11.110 1.180 ;
        RECT  10.510 0.300 10.710 1.180 ;
        RECT  9.220 0.300 10.710 0.460 ;
        RECT  8.160 0.500 9.390 0.870 ;
        RECT  9.220 0.300 9.390 0.870 ;
        RECT  8.160 0.300 8.320 0.870 ;
        RECT  7.300 0.300 8.320 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.350 1.840 13.620 2.540 ;
        RECT  12.270 2.080 12.550 2.540 ;
        RECT  10.020 2.080 10.300 2.540 ;
        RECT  8.600 1.860 8.880 2.540 ;
        RECT  4.780 1.760 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.350 -0.140 13.620 0.560 ;
        RECT  12.270 -0.140 12.550 0.520 ;
        RECT  11.110 -0.140 11.390 0.660 ;
        RECT  8.640 -0.140 8.920 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.100 1.540 0.380 1.920 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.750 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.600 ;
        RECT  4.200 1.440 5.330 1.600 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  5.170 1.440 5.330 2.020 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  5.860 0.620 6.200 1.280 ;
        RECT  4.520 1.120 6.200 1.280 ;
        RECT  5.490 1.120 5.710 1.960 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 6.540 0.460 ;
        RECT  1.150 0.330 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.380 0.300 6.540 1.330 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.220 1.440 2.070 1.600 ;
        RECT  6.700 0.950 7.560 1.230 ;
        RECT  6.700 0.560 6.860 1.960 ;
        RECT  6.070 1.640 6.860 1.960 ;
        RECT  11.300 1.000 11.850 1.160 ;
        RECT  8.160 1.100 10.350 1.320 ;
        RECT  10.070 0.620 10.350 1.600 ;
        RECT  9.360 1.100 10.350 1.600 ;
        RECT  11.300 1.000 11.460 1.600 ;
        RECT  9.360 1.370 11.460 1.600 ;
        RECT  12.570 1.050 13.190 1.270 ;
        RECT  7.720 0.620 8.000 1.960 ;
        RECT  7.020 1.520 8.000 1.960 ;
        RECT  7.020 1.540 9.200 1.700 ;
        RECT  9.040 1.540 9.200 1.920 ;
        RECT  12.570 1.050 12.730 1.920 ;
        RECT  9.040 1.760 12.730 1.920 ;
        RECT  7.020 1.540 8.200 1.960 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.760 2.400 ;
        RECT  9.120 1.080 9.880 2.400 ;
        RECT  10.530 1.080 12.720 2.400 ;
        RECT  0.000 1.140 5.900 2.400 ;
        RECT  7.910 1.140 14.000 2.400 ;
        RECT  0.000 1.260 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.760 0.000 9.120 1.140 ;
        RECT  9.880 0.000 10.530 1.140 ;
        RECT  12.720 0.000 14.000 1.140 ;
        RECT  5.900 0.000 7.910 1.260 ;
    END
END DFRM4HM

MACRO DFRM2HM
    CLASS CORE ;
    FOREIGN DFRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.484  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.210 1.100 0.410 1.300 ;
        LAYER ME2 ;
        RECT  0.100 0.900 0.430 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.020 0.570 1.360 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.900 0.380 11.260 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.080 0.380 12.300 2.100 ;
        RECT  12.020 0.380 12.300 0.700 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.160 0.500 9.220 0.870 ;
        RECT  8.160 0.300 8.320 0.870 ;
        RECT  7.300 0.300 8.320 0.460 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  11.460 2.080 11.740 2.540 ;
        RECT  10.020 2.080 10.300 2.540 ;
        RECT  8.600 1.860 8.880 2.540 ;
        RECT  4.780 1.760 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  11.460 -0.140 11.740 0.520 ;
        RECT  10.480 -0.140 10.680 0.660 ;
        RECT  8.640 -0.140 8.920 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.100 1.540 0.380 1.920 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.750 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.600 ;
        RECT  4.200 1.440 5.330 1.600 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  5.170 1.440 5.330 2.020 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  5.860 0.620 6.200 1.280 ;
        RECT  4.520 1.120 6.200 1.280 ;
        RECT  5.490 1.120 5.710 1.960 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 6.540 0.460 ;
        RECT  1.150 0.310 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.380 0.300 6.540 1.330 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.220 1.440 2.070 1.600 ;
        RECT  6.700 0.950 7.560 1.230 ;
        RECT  6.700 0.560 6.860 1.960 ;
        RECT  6.070 1.640 6.860 1.960 ;
        RECT  10.000 0.400 10.200 1.260 ;
        RECT  10.000 1.000 10.710 1.260 ;
        RECT  8.160 1.100 10.710 1.260 ;
        RECT  9.390 1.100 9.690 1.600 ;
        RECT  7.720 0.620 8.000 1.960 ;
        RECT  7.020 1.520 8.000 1.960 ;
        RECT  7.020 1.540 9.200 1.700 ;
        RECT  9.040 1.540 9.200 1.920 ;
        RECT  11.730 0.950 11.890 1.920 ;
        RECT  9.040 1.760 11.890 1.920 ;
        RECT  7.020 1.540 8.200 1.960 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.760 2.400 ;
        RECT  9.120 1.080 11.440 2.400 ;
        RECT  0.000 1.140 5.900 2.400 ;
        RECT  7.890 1.140 12.400 2.400 ;
        RECT  0.000 1.260 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.760 0.000 9.120 1.140 ;
        RECT  11.440 0.000 12.400 1.140 ;
        RECT  5.900 0.000 7.890 1.260 ;
    END
END DFRM2HM

MACRO DFRM1HM
    CLASS CORE ;
    FOREIGN DFRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.900 0.380 11.260 1.600 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.370 1.100 2.570 1.300 ;
        LAYER ME2 ;
        RECT  2.370 0.900 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.260 1.010 2.570 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.068  LAYER ME1  ;
        ANTENNAGATEAREA 0.068  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.158  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.220 1.080 0.420 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.420 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.020 0.570 1.360 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.080 0.380 12.300 2.100 ;
        RECT  12.020 0.380 12.300 0.700 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.160 0.500 9.220 0.870 ;
        RECT  8.160 0.300 8.320 0.870 ;
        RECT  7.300 0.300 8.320 0.460 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  11.460 2.080 11.740 2.540 ;
        RECT  10.020 2.080 10.300 2.540 ;
        RECT  8.600 1.860 8.880 2.540 ;
        RECT  4.780 1.760 4.940 2.540 ;
        RECT  3.760 1.500 4.040 2.540 ;
        RECT  1.600 2.080 1.880 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  11.460 -0.140 11.740 0.520 ;
        RECT  10.480 -0.140 10.680 0.660 ;
        RECT  8.640 -0.140 8.920 0.320 ;
        RECT  5.160 -0.140 5.380 0.600 ;
        RECT  4.170 -0.140 4.450 0.320 ;
        RECT  1.630 -0.140 1.910 0.380 ;
        RECT  0.630 -0.140 0.910 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 0.380 0.860 ;
        RECT  0.100 0.700 0.910 0.860 ;
        RECT  0.730 0.700 0.910 1.260 ;
        RECT  0.730 1.040 1.570 1.260 ;
        RECT  0.100 1.540 0.380 1.920 ;
        RECT  0.730 0.700 0.890 1.920 ;
        RECT  0.100 1.750 0.890 1.920 ;
        RECT  0.100 1.760 2.200 1.920 ;
        RECT  2.040 1.760 2.200 2.100 ;
        RECT  2.040 1.940 3.220 2.100 ;
        RECT  2.610 0.620 2.890 0.840 ;
        RECT  2.730 1.180 4.360 1.340 ;
        RECT  4.200 1.180 4.360 1.600 ;
        RECT  4.200 1.440 5.330 1.600 ;
        RECT  2.730 0.620 2.890 1.780 ;
        RECT  2.510 1.560 2.890 1.780 ;
        RECT  5.170 1.440 5.330 2.020 ;
        RECT  3.430 0.860 4.680 1.020 ;
        RECT  4.520 0.860 4.680 1.280 ;
        RECT  5.860 0.620 6.200 1.280 ;
        RECT  4.520 1.120 6.200 1.280 ;
        RECT  5.490 1.120 5.710 1.920 ;
        RECT  2.070 0.300 3.210 0.460 ;
        RECT  5.540 0.300 6.540 0.460 ;
        RECT  1.150 0.310 1.430 0.700 ;
        RECT  3.050 0.300 3.210 1.020 ;
        RECT  2.070 0.300 2.250 0.700 ;
        RECT  1.150 0.540 2.250 0.700 ;
        RECT  3.050 0.540 5.000 0.700 ;
        RECT  4.840 0.540 5.000 0.920 ;
        RECT  5.540 0.300 5.700 0.920 ;
        RECT  4.840 0.760 5.700 0.920 ;
        RECT  3.050 0.540 3.250 1.020 ;
        RECT  6.380 0.300 6.540 1.330 ;
        RECT  1.910 0.540 2.070 1.600 ;
        RECT  1.220 1.440 2.070 1.600 ;
        RECT  6.700 0.950 7.560 1.230 ;
        RECT  6.700 0.560 6.860 1.920 ;
        RECT  6.070 1.640 6.860 1.920 ;
        RECT  10.000 0.340 10.200 1.260 ;
        RECT  10.000 1.000 10.720 1.260 ;
        RECT  8.160 1.100 10.720 1.260 ;
        RECT  9.390 1.100 9.690 1.600 ;
        RECT  7.720 0.620 8.000 1.960 ;
        RECT  7.720 1.540 9.200 1.700 ;
        RECT  9.040 1.540 9.200 1.920 ;
        RECT  11.730 0.950 11.890 1.920 ;
        RECT  9.040 1.760 11.890 1.920 ;
        RECT  7.020 1.680 8.200 1.960 ;
        LAYER VTPH ;
        RECT  0.930 1.080 1.760 2.400 ;
        RECT  9.120 1.080 11.440 2.400 ;
        RECT  0.000 1.140 5.900 2.400 ;
        RECT  7.640 1.140 12.400 2.400 ;
        RECT  0.000 1.260 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.080 ;
        RECT  0.000 0.000 0.930 1.140 ;
        RECT  1.760 0.000 9.120 1.140 ;
        RECT  11.440 0.000 12.400 1.140 ;
        RECT  5.900 0.000 7.640 1.260 ;
    END
END DFRM1HM

MACRO DFQZRM8HM
    CLASS CORE ;
    FOREIGN DFQZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.460 0.900 11.750 2.100 ;
        RECT  11.470 0.380 11.750 2.100 ;
        RECT  10.550 0.900 11.750 1.200 ;
        RECT  10.430 1.470 10.710 2.100 ;
        RECT  10.550 0.380 10.710 2.100 ;
        RECT  10.430 0.380 10.710 0.780 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  12.030 1.470 12.230 2.540 ;
        RECT  10.990 1.470 11.190 2.540 ;
        RECT  9.950 1.470 10.150 2.540 ;
        RECT  8.910 1.470 9.110 2.540 ;
        RECT  7.610 1.970 7.770 2.540 ;
        RECT  4.790 2.080 5.070 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  11.990 -0.140 12.270 0.620 ;
        RECT  10.990 -0.140 11.190 0.680 ;
        RECT  9.950 -0.140 10.150 0.700 ;
        RECT  8.910 -0.140 9.110 0.630 ;
        RECT  7.520 -0.140 7.800 0.320 ;
        RECT  4.790 -0.140 5.070 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.710 0.920 5.330 1.080 ;
        RECT  3.710 0.640 3.990 1.780 ;
        RECT  4.370 1.240 5.750 1.400 ;
        RECT  5.550 0.620 5.750 1.780 ;
        RECT  0.140 0.400 0.340 0.680 ;
        RECT  0.140 0.520 1.180 0.680 ;
        RECT  0.940 0.520 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.250 1.760 5.390 1.920 ;
        RECT  1.020 0.520 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.230 1.760 5.390 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.250 1.760 4.410 2.100 ;
        RECT  2.780 1.940 4.410 2.100 ;
        RECT  5.950 1.200 6.110 2.100 ;
        RECT  5.230 1.940 6.110 2.100 ;
        RECT  3.340 0.300 4.410 0.460 ;
        RECT  5.230 0.300 6.750 0.460 ;
        RECT  4.250 0.300 4.410 0.640 ;
        RECT  5.230 0.300 5.390 0.640 ;
        RECT  4.250 0.480 5.390 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.590 0.300 6.750 1.650 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.970 0.480 8.430 0.640 ;
        RECT  6.970 1.320 8.430 1.480 ;
        RECT  6.970 0.480 7.130 1.780 ;
        RECT  8.270 1.320 8.430 1.780 ;
        RECT  6.070 0.640 6.430 0.800 ;
        RECT  8.590 1.120 9.190 1.280 ;
        RECT  7.290 1.640 8.110 1.800 ;
        RECT  6.270 0.640 6.430 2.100 ;
        RECT  7.950 1.640 8.110 2.100 ;
        RECT  7.290 1.640 7.450 2.100 ;
        RECT  6.270 1.940 7.450 2.100 ;
        RECT  8.590 1.120 8.750 2.100 ;
        RECT  7.950 1.940 8.750 2.100 ;
        RECT  7.760 0.800 9.690 0.960 ;
        RECT  9.350 0.430 9.690 1.280 ;
        RECT  7.760 0.800 8.050 1.160 ;
        RECT  9.350 1.000 10.330 1.280 ;
        RECT  9.350 0.430 9.670 2.100 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  4.130 1.140 5.090 2.400 ;
        RECT  0.000 1.160 5.090 2.400 ;
        RECT  6.530 1.140 12.400 2.400 ;
        RECT  0.000 1.200 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 12.400 1.140 ;
        RECT  3.400 0.000 4.130 1.160 ;
        RECT  5.090 0.000 6.530 1.200 ;
    END
END DFQZRM8HM

MACRO DFQZRM4HM
    CLASS CORE ;
    FOREIGN DFQZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.645  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.250 0.470 8.410 1.760 ;
        RECT  8.100 0.470 8.410 1.160 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.930 1.480 10.130 2.540 ;
        RECT  8.890 1.840 9.090 2.540 ;
        RECT  7.610 1.760 7.770 2.540 ;
        RECT  4.790 2.080 5.070 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.950 -0.140 10.110 0.760 ;
        RECT  8.710 -0.140 8.990 0.590 ;
        RECT  7.530 -0.140 7.730 0.680 ;
        RECT  4.790 -0.140 5.070 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.710 0.920 5.330 1.080 ;
        RECT  3.710 0.640 3.990 1.780 ;
        RECT  4.370 1.240 5.750 1.400 ;
        RECT  5.550 0.620 5.750 1.780 ;
        RECT  0.100 0.480 1.180 0.680 ;
        RECT  0.940 0.480 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.250 1.760 5.390 1.920 ;
        RECT  1.020 0.480 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.230 1.760 5.390 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.250 1.760 4.410 2.100 ;
        RECT  2.780 1.940 4.410 2.100 ;
        RECT  5.950 1.200 6.110 2.100 ;
        RECT  5.230 1.940 6.110 2.100 ;
        RECT  3.340 0.300 4.410 0.460 ;
        RECT  5.230 0.300 6.750 0.460 ;
        RECT  4.250 0.300 4.410 0.640 ;
        RECT  5.230 0.300 5.390 0.640 ;
        RECT  4.250 0.480 5.390 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  6.590 0.300 6.750 1.680 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.970 0.380 7.130 1.780 ;
        RECT  6.070 0.640 6.430 0.800 ;
        RECT  8.890 1.120 9.330 1.280 ;
        RECT  7.290 1.390 8.090 1.550 ;
        RECT  8.890 1.120 9.050 1.680 ;
        RECT  8.570 1.520 9.050 1.680 ;
        RECT  6.270 0.640 6.430 2.100 ;
        RECT  7.930 1.390 8.090 2.100 ;
        RECT  7.290 1.390 7.450 2.100 ;
        RECT  6.270 1.940 7.450 2.100 ;
        RECT  8.570 1.520 8.730 2.100 ;
        RECT  7.930 1.940 8.730 2.100 ;
        RECT  9.360 0.390 9.670 0.960 ;
        RECT  8.570 0.800 9.670 0.960 ;
        RECT  8.570 0.800 8.730 1.360 ;
        RECT  9.490 0.390 9.670 2.100 ;
        RECT  9.370 1.480 9.670 2.100 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  0.000 1.160 5.090 2.400 ;
        RECT  6.700 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 10.400 1.140 ;
        RECT  3.400 0.000 6.700 1.160 ;
        RECT  5.090 0.000 6.700 1.200 ;
    END
END DFQZRM4HM

MACRO DFQZRM2HM
    CLASS CORE ;
    FOREIGN DFQZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.418  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.240 0.460 8.400 1.760 ;
        RECT  8.040 1.300 8.400 1.500 ;
        RECT  8.120 0.460 8.400 1.500 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.220 1.630 9.420 2.540 ;
        RECT  7.560 2.020 7.760 2.540 ;
        RECT  4.740 2.080 5.020 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.240 -0.140 9.400 0.840 ;
        RECT  7.380 -0.140 7.660 0.670 ;
        RECT  4.740 -0.140 5.020 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.660 0.920 5.280 1.080 ;
        RECT  3.660 0.640 3.940 1.780 ;
        RECT  4.320 1.240 5.700 1.400 ;
        RECT  5.500 0.620 5.700 1.780 ;
        RECT  0.100 0.480 1.180 0.680 ;
        RECT  0.940 0.480 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.200 1.760 5.340 1.920 ;
        RECT  1.020 0.480 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.180 1.760 5.340 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.200 1.760 4.360 2.100 ;
        RECT  2.780 1.940 4.360 2.100 ;
        RECT  5.900 1.200 6.060 2.100 ;
        RECT  5.180 1.940 6.060 2.100 ;
        RECT  3.340 0.300 4.360 0.460 ;
        RECT  5.180 0.300 6.700 0.460 ;
        RECT  4.200 0.300 4.360 0.640 ;
        RECT  5.180 0.300 5.340 0.640 ;
        RECT  4.200 0.480 5.340 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.540 0.300 6.700 1.620 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.910 0.360 7.080 1.780 ;
        RECT  6.020 0.640 6.380 0.800 ;
        RECT  7.240 1.700 8.080 1.860 ;
        RECT  6.220 0.640 6.380 2.100 ;
        RECT  7.920 1.700 8.080 2.100 ;
        RECT  7.240 1.700 7.400 2.100 ;
        RECT  6.220 1.940 7.400 2.100 ;
        RECT  7.920 1.940 8.640 2.100 ;
        RECT  8.580 1.040 8.940 1.320 ;
        RECT  8.660 0.460 8.940 1.660 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  0.000 1.160 5.040 2.400 ;
        RECT  6.570 1.140 9.600 2.400 ;
        RECT  0.000 1.200 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 9.600 1.140 ;
        RECT  3.400 0.000 6.570 1.160 ;
        RECT  5.040 0.000 6.570 1.200 ;
    END
END DFQZRM2HM

MACRO DFQZRM1HM
    CLASS CORE ;
    FOREIGN DFQZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.840 2.800 1.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.314  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.240 0.570 8.400 1.760 ;
        RECT  8.040 1.300 8.400 1.500 ;
        RECT  8.120 0.570 8.400 1.500 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.220 1.530 9.420 2.540 ;
        RECT  7.560 2.020 7.760 2.540 ;
        RECT  4.740 2.080 5.020 2.540 ;
        RECT  2.340 2.080 2.620 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.240 -0.140 9.400 0.840 ;
        RECT  7.380 -0.140 7.660 0.670 ;
        RECT  4.740 -0.140 5.020 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.380 3.180 1.600 ;
        RECT  1.740 1.440 3.180 1.600 ;
        RECT  3.660 0.920 5.280 1.080 ;
        RECT  3.660 0.640 3.940 1.780 ;
        RECT  4.320 1.240 5.700 1.400 ;
        RECT  5.500 0.620 5.700 1.780 ;
        RECT  0.100 0.480 1.180 0.680 ;
        RECT  0.940 0.480 1.180 1.680 ;
        RECT  0.140 1.520 1.180 1.680 ;
        RECT  1.780 1.760 2.940 1.920 ;
        RECT  4.200 1.760 5.340 1.920 ;
        RECT  1.020 0.480 1.180 2.100 ;
        RECT  2.780 1.760 2.940 2.100 ;
        RECT  5.180 1.760 5.340 2.100 ;
        RECT  0.140 1.520 0.340 2.040 ;
        RECT  1.780 1.760 1.940 2.100 ;
        RECT  1.020 1.940 1.940 2.100 ;
        RECT  4.200 1.760 4.360 2.100 ;
        RECT  2.780 1.940 4.360 2.100 ;
        RECT  5.900 1.200 6.060 2.100 ;
        RECT  5.180 1.940 6.060 2.100 ;
        RECT  3.340 0.300 4.360 0.460 ;
        RECT  5.180 0.300 6.700 0.460 ;
        RECT  4.200 0.300 4.360 0.640 ;
        RECT  5.180 0.300 5.340 0.640 ;
        RECT  4.200 0.480 5.340 0.640 ;
        RECT  1.340 0.480 3.500 0.680 ;
        RECT  6.540 0.300 6.700 1.590 ;
        RECT  3.340 0.300 3.500 1.660 ;
        RECT  1.340 0.480 1.540 1.760 ;
        RECT  6.910 0.360 7.080 1.780 ;
        RECT  6.020 0.620 6.380 0.780 ;
        RECT  7.240 1.700 8.080 1.860 ;
        RECT  6.220 0.620 6.380 2.100 ;
        RECT  7.920 1.700 8.080 2.100 ;
        RECT  7.240 1.700 7.400 2.100 ;
        RECT  6.220 1.940 7.400 2.100 ;
        RECT  7.920 1.940 8.640 2.100 ;
        RECT  8.580 1.040 8.940 1.320 ;
        RECT  8.660 0.570 8.940 1.660 ;
        LAYER VTPH ;
        RECT  1.540 1.080 3.400 2.400 ;
        RECT  0.000 1.140 3.400 2.400 ;
        RECT  0.000 1.160 5.040 2.400 ;
        RECT  6.570 1.140 9.600 2.400 ;
        RECT  0.000 1.200 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.080 ;
        RECT  0.000 0.000 1.540 1.140 ;
        RECT  3.400 0.000 9.600 1.140 ;
        RECT  3.400 0.000 6.570 1.160 ;
        RECT  5.040 0.000 6.570 1.200 ;
    END
END DFQZRM1HM

MACRO DFQSM8HM
    CLASS CORE ;
    FOREIGN DFQSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.154  LAYER ME1  ;
        ANTENNAGATEAREA 0.154  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 16.318  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.020 7.100 1.220 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.800 1.020 7.410 1.220 ;
        RECT  7.250 0.300 7.410 1.220 ;
        RECT  5.350 0.300 7.410 0.460 ;
        RECT  4.800 1.020 5.510 1.300 ;
        RECT  5.350 0.300 5.510 1.300 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        ANTENNAGATEAREA 0.127  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.352  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.140 2.700 1.340 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.410 1.030 2.800 1.460 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.470 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.720 1.000 11.100 1.300 ;
        RECT  10.740 0.800 11.100 1.300 ;
        RECT  10.740 0.430 10.940 2.080 ;
        RECT  9.720 1.000 9.920 2.080 ;
        RECT  9.720 0.390 9.880 2.080 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.260 1.470 11.460 2.540 ;
        RECT  10.220 1.480 10.420 2.540 ;
        RECT  9.180 1.480 9.380 2.540 ;
        RECT  8.140 1.840 8.340 2.540 ;
        RECT  4.790 1.860 5.070 2.540 ;
        RECT  3.670 1.860 3.950 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.260 -0.140 11.460 0.710 ;
        RECT  10.220 -0.140 10.420 0.710 ;
        RECT  9.180 -0.140 9.380 0.710 ;
        RECT  7.930 -0.140 8.130 0.560 ;
        RECT  3.710 -0.140 3.910 0.380 ;
        RECT  1.750 -0.140 2.050 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.440 0.920 0.640 ;
        RECT  0.740 1.010 1.640 1.210 ;
        RECT  0.740 0.440 0.920 1.920 ;
        RECT  0.100 1.720 0.920 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.290 2.100 ;
        RECT  2.730 0.640 3.120 0.840 ;
        RECT  2.960 0.640 3.120 1.780 ;
        RECT  2.960 0.900 4.120 1.060 ;
        RECT  3.920 0.900 4.120 1.260 ;
        RECT  2.960 0.900 3.150 1.780 ;
        RECT  2.500 1.620 3.150 1.780 ;
        RECT  2.330 0.300 3.510 0.460 ;
        RECT  4.150 0.300 5.190 0.460 ;
        RECT  4.910 0.300 5.190 0.500 ;
        RECT  3.350 0.300 3.510 0.720 ;
        RECT  4.150 0.300 4.310 0.720 ;
        RECT  3.350 0.550 4.310 0.720 ;
        RECT  1.150 0.530 2.510 0.760 ;
        RECT  2.330 0.300 2.510 0.790 ;
        RECT  1.930 0.530 2.510 0.790 ;
        RECT  1.930 0.530 2.090 1.600 ;
        RECT  1.110 1.400 2.090 1.600 ;
        RECT  4.470 0.640 4.830 0.840 ;
        RECT  3.410 1.240 3.610 1.700 ;
        RECT  4.470 0.640 4.640 1.700 ;
        RECT  3.410 1.540 5.510 1.700 ;
        RECT  5.310 1.540 5.510 1.850 ;
        RECT  6.210 0.620 7.090 0.840 ;
        RECT  6.210 0.620 6.370 1.780 ;
        RECT  6.210 1.500 7.660 1.660 ;
        RECT  6.210 1.500 6.680 1.780 ;
        RECT  8.100 1.050 8.300 1.680 ;
        RECT  7.820 1.520 8.300 1.680 ;
        RECT  5.670 0.640 5.870 1.720 ;
        RECT  5.860 1.520 6.020 2.100 ;
        RECT  7.820 1.520 7.980 2.100 ;
        RECT  5.860 1.940 7.980 2.100 ;
        RECT  7.570 0.730 8.860 0.890 ;
        RECT  8.660 1.000 9.560 1.200 ;
        RECT  7.570 0.730 7.730 1.280 ;
        RECT  8.660 0.430 8.860 2.080 ;
        LAYER VTPH ;
        RECT  0.530 1.080 2.100 2.400 ;
        RECT  0.000 1.140 2.100 2.400 ;
        RECT  3.570 1.160 5.310 2.400 ;
        RECT  0.000 1.200 5.310 2.400 ;
        RECT  6.700 1.140 11.600 2.400 ;
        RECT  0.000 1.240 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.080 ;
        RECT  0.000 0.000 0.530 1.140 ;
        RECT  2.100 0.000 11.600 1.140 ;
        RECT  2.100 0.000 6.700 1.160 ;
        RECT  2.100 0.000 3.570 1.200 ;
        RECT  5.310 0.000 6.700 1.240 ;
    END
END DFQSM8HM

MACRO DFQSM4HM
    CLASS CORE ;
    FOREIGN DFQSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 17.595  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.020 7.100 1.220 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.800 1.020 7.300 1.220 ;
        RECT  7.140 0.300 7.300 1.220 ;
        RECT  5.240 0.300 7.300 0.460 ;
        RECT  4.690 1.020 5.400 1.300 ;
        RECT  5.240 0.300 5.400 1.300 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.470 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.190 2.580 1.390 ;
        RECT  2.100 1.190 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.490 0.840 9.900 1.160 ;
        RECT  9.490 0.390 9.700 2.080 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  10.010 1.480 10.210 2.540 ;
        RECT  8.970 1.480 9.170 2.540 ;
        RECT  7.930 1.840 8.130 2.540 ;
        RECT  4.680 1.860 4.960 2.540 ;
        RECT  3.560 1.860 3.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  10.010 -0.140 10.210 0.710 ;
        RECT  8.970 -0.140 9.170 0.710 ;
        RECT  7.660 -0.140 7.860 0.560 ;
        RECT  3.460 -0.140 3.660 0.380 ;
        RECT  1.660 -0.140 1.860 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.530 0.920 0.730 ;
        RECT  0.740 0.920 1.330 1.120 ;
        RECT  0.740 0.530 0.920 1.920 ;
        RECT  0.100 1.720 0.920 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.180 2.100 ;
        RECT  2.560 0.680 2.920 0.840 ;
        RECT  2.760 0.900 4.010 1.060 ;
        RECT  3.810 0.900 4.010 1.260 ;
        RECT  2.760 0.680 2.920 1.780 ;
        RECT  2.480 1.580 2.920 1.780 ;
        RECT  2.020 0.300 3.260 0.460 ;
        RECT  4.040 0.300 5.080 0.460 ;
        RECT  4.800 0.300 5.080 0.500 ;
        RECT  3.100 0.300 3.260 0.720 ;
        RECT  4.040 0.300 4.200 0.720 ;
        RECT  3.100 0.550 4.200 0.720 ;
        RECT  2.020 0.300 2.200 0.740 ;
        RECT  1.140 0.540 2.200 0.740 ;
        RECT  1.590 0.540 1.790 1.600 ;
        RECT  1.100 1.400 1.790 1.600 ;
        RECT  4.360 0.640 4.720 0.840 ;
        RECT  3.290 1.240 3.490 1.700 ;
        RECT  4.360 0.640 4.530 1.700 ;
        RECT  3.290 1.540 5.400 1.700 ;
        RECT  5.200 1.540 5.400 1.850 ;
        RECT  6.100 0.620 6.980 0.840 ;
        RECT  6.100 0.620 6.260 1.780 ;
        RECT  6.100 1.580 7.450 1.780 ;
        RECT  8.090 1.050 8.290 1.680 ;
        RECT  7.610 1.520 8.290 1.680 ;
        RECT  5.560 0.640 5.760 1.720 ;
        RECT  5.750 1.520 5.910 2.100 ;
        RECT  7.610 1.520 7.770 2.100 ;
        RECT  5.750 1.940 7.770 2.100 ;
        RECT  7.460 0.730 8.650 0.890 ;
        RECT  8.450 0.960 9.290 1.240 ;
        RECT  7.460 0.730 7.620 1.280 ;
        RECT  8.450 0.430 8.650 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.080 1.750 2.400 ;
        RECT  3.570 1.160 5.200 2.400 ;
        RECT  0.000 1.200 5.200 2.400 ;
        RECT  6.590 1.140 10.400 2.400 ;
        RECT  0.000 1.240 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  1.750 0.000 10.400 1.140 ;
        RECT  1.750 0.000 6.590 1.160 ;
        RECT  1.750 0.000 3.570 1.200 ;
        RECT  5.200 0.000 6.590 1.240 ;
    END
END DFQSM4HM

MACRO DFQSM2HM
    CLASS CORE ;
    FOREIGN DFQSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.139  LAYER ME1  ;
        ANTENNAGATEAREA 0.139  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 17.595  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.020 7.100 1.220 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.800 1.020 7.300 1.220 ;
        RECT  7.140 0.300 7.300 1.220 ;
        RECT  5.240 0.300 7.300 0.460 ;
        RECT  4.690 1.020 5.400 1.300 ;
        RECT  5.240 0.300 5.400 1.300 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.470 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.190 2.580 1.390 ;
        RECT  2.100 1.190 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.300 0.390 9.590 2.080 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  8.890 1.840 9.090 2.540 ;
        RECT  7.930 1.840 8.130 2.540 ;
        RECT  4.680 1.860 4.960 2.540 ;
        RECT  3.560 1.860 3.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  8.890 -0.140 9.090 0.710 ;
        RECT  7.750 -0.140 7.950 0.560 ;
        RECT  3.460 -0.140 3.660 0.380 ;
        RECT  1.660 -0.140 1.860 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.530 0.920 0.730 ;
        RECT  0.740 0.920 1.330 1.120 ;
        RECT  0.740 0.530 0.920 1.920 ;
        RECT  0.100 1.720 0.920 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.180 2.100 ;
        RECT  2.560 0.680 2.920 0.840 ;
        RECT  2.760 0.900 4.010 1.060 ;
        RECT  3.810 0.900 4.010 1.260 ;
        RECT  2.760 0.680 2.920 1.780 ;
        RECT  2.480 1.580 2.920 1.780 ;
        RECT  2.020 0.300 3.260 0.460 ;
        RECT  4.040 0.300 5.080 0.460 ;
        RECT  4.800 0.300 5.080 0.500 ;
        RECT  3.100 0.300 3.260 0.720 ;
        RECT  4.040 0.300 4.200 0.720 ;
        RECT  3.100 0.550 4.200 0.720 ;
        RECT  2.020 0.300 2.200 0.740 ;
        RECT  1.140 0.540 2.200 0.740 ;
        RECT  1.590 0.540 1.790 1.600 ;
        RECT  1.100 1.400 1.790 1.600 ;
        RECT  4.360 0.640 4.720 0.840 ;
        RECT  3.290 1.240 3.490 1.700 ;
        RECT  4.360 0.640 4.530 1.700 ;
        RECT  3.290 1.540 5.400 1.700 ;
        RECT  5.200 1.540 5.400 1.850 ;
        RECT  6.100 0.620 6.980 0.840 ;
        RECT  6.100 0.620 6.260 1.780 ;
        RECT  6.100 1.580 7.450 1.780 ;
        RECT  7.940 1.050 8.140 1.680 ;
        RECT  7.610 1.520 8.140 1.680 ;
        RECT  5.560 0.640 5.760 1.720 ;
        RECT  5.750 1.520 5.910 2.100 ;
        RECT  7.610 1.520 7.770 2.100 ;
        RECT  5.750 1.940 7.770 2.100 ;
        RECT  8.270 0.430 8.470 0.890 ;
        RECT  7.460 0.730 8.470 0.890 ;
        RECT  8.300 0.430 8.470 1.200 ;
        RECT  8.300 1.000 9.050 1.200 ;
        RECT  7.460 0.730 7.620 1.280 ;
        RECT  8.450 1.000 8.650 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.080 1.750 2.400 ;
        RECT  3.570 1.160 5.200 2.400 ;
        RECT  0.000 1.200 5.200 2.400 ;
        RECT  6.590 1.140 10.000 2.400 ;
        RECT  0.000 1.240 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.080 ;
        RECT  1.750 0.000 10.000 1.140 ;
        RECT  1.750 0.000 6.590 1.160 ;
        RECT  1.750 0.000 3.570 1.200 ;
        RECT  5.200 0.000 6.590 1.240 ;
    END
END DFQSM2HM

MACRO DFQSM1HM
    CLASS CORE ;
    FOREIGN DFQSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 20.616  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.900 1.020 7.100 1.220 ;
        LAYER ME2 ;
        RECT  6.900 0.840 7.100 1.560 ;
        LAYER ME1 ;
        RECT  6.800 1.020 7.300 1.220 ;
        RECT  7.140 0.300 7.300 1.220 ;
        RECT  5.240 0.300 7.300 0.460 ;
        RECT  4.690 1.020 5.400 1.300 ;
        RECT  5.240 0.300 5.400 1.300 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.470 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.190 2.580 1.390 ;
        RECT  2.100 1.190 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.490 0.820 9.900 1.220 ;
        RECT  9.490 0.390 9.700 2.080 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  8.970 1.840 9.170 2.540 ;
        RECT  7.930 1.840 8.130 2.540 ;
        RECT  4.680 1.860 4.960 2.540 ;
        RECT  3.560 1.860 3.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  8.970 -0.140 9.170 0.670 ;
        RECT  7.750 -0.140 7.950 0.560 ;
        RECT  3.460 -0.140 3.660 0.380 ;
        RECT  1.660 -0.140 1.860 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.540 0.920 0.740 ;
        RECT  0.740 0.920 1.330 1.120 ;
        RECT  0.740 0.540 0.920 1.920 ;
        RECT  0.100 1.720 0.920 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.180 2.100 ;
        RECT  2.560 0.680 2.920 0.840 ;
        RECT  2.760 0.900 4.010 1.060 ;
        RECT  3.810 0.900 4.010 1.260 ;
        RECT  2.760 0.680 2.920 1.780 ;
        RECT  2.480 1.580 2.920 1.780 ;
        RECT  2.020 0.300 3.260 0.460 ;
        RECT  4.040 0.300 5.080 0.460 ;
        RECT  4.800 0.300 5.080 0.500 ;
        RECT  3.100 0.300 3.260 0.720 ;
        RECT  4.040 0.300 4.200 0.720 ;
        RECT  3.100 0.550 4.200 0.720 ;
        RECT  2.020 0.300 2.200 0.740 ;
        RECT  1.140 0.540 2.200 0.740 ;
        RECT  1.590 0.540 1.790 1.600 ;
        RECT  1.100 1.400 1.790 1.600 ;
        RECT  4.360 0.640 4.720 0.840 ;
        RECT  3.290 1.240 3.490 1.700 ;
        RECT  4.360 0.640 4.530 1.700 ;
        RECT  3.290 1.540 5.400 1.700 ;
        RECT  5.200 1.540 5.400 1.840 ;
        RECT  6.100 0.620 6.980 0.840 ;
        RECT  6.100 0.620 6.260 1.780 ;
        RECT  6.100 1.580 7.450 1.780 ;
        RECT  7.940 1.050 8.140 1.680 ;
        RECT  7.610 1.520 8.140 1.680 ;
        RECT  5.560 0.620 5.760 1.720 ;
        RECT  5.750 1.520 5.910 2.100 ;
        RECT  7.610 1.520 7.770 2.100 ;
        RECT  5.750 1.940 7.770 2.100 ;
        RECT  7.460 0.730 8.690 0.890 ;
        RECT  8.490 1.000 9.180 1.200 ;
        RECT  7.460 0.730 7.620 1.280 ;
        RECT  8.490 0.350 8.690 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.080 1.750 2.400 ;
        RECT  3.570 1.180 5.200 2.400 ;
        RECT  0.000 1.200 5.200 2.400 ;
        RECT  6.590 1.140 10.000 2.400 ;
        RECT  0.000 1.240 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.080 ;
        RECT  1.750 0.000 10.000 1.140 ;
        RECT  1.750 0.000 6.590 1.180 ;
        RECT  1.750 0.000 3.570 1.200 ;
        RECT  5.200 0.000 6.590 1.240 ;
    END
END DFQSM1HM

MACRO DFQRSM8HM
    CLASS CORE ;
    FOREIGN DFQRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 0.320 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.110 2.640 1.310 ;
        RECT  2.100 1.110 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 3.940 1.900 4.420 ;
        RECT  0.500 3.060 1.900 3.260 ;
        RECT  1.700 2.980 1.900 3.260 ;
        RECT  0.500 3.940 1.900 4.140 ;
        RECT  0.500 2.720 0.860 4.420 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.293  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 3.610 4.240 3.810 ;
        RECT  2.500 3.240 2.750 3.810 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 3.640 5.100 4.260 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  3.220 3.080 3.580 3.280 ;
        RECT  3.220 2.260 3.380 3.280 ;
        RECT  2.220 2.260 2.500 2.680 ;
        RECT  1.660 2.140 1.940 2.540 ;
        RECT  1.140 2.260 1.420 2.900 ;
        RECT  0.660 2.140 0.940 2.540 ;
        RECT  0.140 2.260 0.340 3.320 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  4.220 -0.140 4.500 0.320 ;
        RECT  1.700 -0.140 1.980 0.550 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 7.200 4.940 ;
        RECT  4.140 4.300 4.420 4.940 ;
        RECT  2.220 4.300 2.500 4.940 ;
        RECT  1.140 4.300 1.420 4.940 ;
        RECT  0.140 4.140 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.300 1.520 4.180 1.760 ;
        RECT  2.180 2.840 3.060 3.040 ;
        RECT  3.820 3.080 4.740 3.280 ;
        RECT  1.120 3.520 2.340 3.720 ;
        RECT  2.180 2.840 2.340 4.140 ;
        RECT  4.580 3.080 4.740 4.140 ;
        RECT  2.180 3.970 4.740 4.140 ;
        RECT  3.340 3.970 3.540 4.360 ;
        RECT  2.520 0.640 2.960 0.800 ;
        RECT  2.800 0.800 4.820 0.960 ;
        RECT  4.660 0.800 4.820 1.380 ;
        RECT  2.800 0.640 2.960 1.760 ;
        RECT  2.500 1.600 2.960 1.760 ;
        RECT  2.140 0.320 3.280 0.480 ;
        RECT  3.120 0.480 5.140 0.640 ;
        RECT  1.260 0.440 1.460 0.870 ;
        RECT  2.140 0.320 2.300 0.870 ;
        RECT  1.260 0.710 2.300 0.870 ;
        RECT  4.980 0.480 5.140 1.210 ;
        RECT  4.980 1.010 5.880 1.210 ;
        RECT  1.420 0.710 1.580 1.660 ;
        RECT  1.180 1.500 1.580 1.660 ;
        RECT  0.140 0.440 0.340 0.860 ;
        RECT  0.140 0.700 0.640 0.860 ;
        RECT  0.480 1.100 1.040 1.300 ;
        RECT  0.480 0.700 0.640 1.980 ;
        RECT  0.140 1.720 0.640 1.980 ;
        RECT  0.140 1.820 2.240 1.980 ;
        RECT  0.140 1.720 0.340 2.000 ;
        RECT  2.090 1.920 6.200 2.080 ;
        RECT  5.300 0.500 5.500 0.780 ;
        RECT  5.300 0.620 6.200 0.780 ;
        RECT  3.480 1.120 4.500 1.280 ;
        RECT  4.340 1.120 4.500 1.700 ;
        RECT  6.040 0.620 6.200 1.700 ;
        RECT  4.340 1.540 6.200 1.700 ;
        RECT  4.940 3.200 6.380 3.360 ;
        RECT  5.340 3.200 6.380 3.420 ;
        RECT  5.340 3.200 5.540 4.480 ;
        RECT  6.420 0.350 6.620 1.760 ;
        RECT  3.600 2.720 6.950 2.880 ;
        RECT  6.790 2.720 6.950 4.480 ;
        RECT  6.100 4.280 6.950 4.480 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.300 3.660 ;
        RECT  3.100 1.140 7.200 3.660 ;
        RECT  0.000 1.200 7.200 3.660 ;
        RECT  4.800 1.140 6.560 3.720 ;
        LAYER VTNH ;
        RECT  0.000 3.660 4.800 4.800 ;
        RECT  6.560 3.660 7.200 4.800 ;
        RECT  0.000 3.720 7.200 4.800 ;
        RECT  0.000 0.000 7.200 1.140 ;
        RECT  2.300 0.000 3.100 1.200 ;
    END
END DFQRSM8HM

MACRO DFQRSM4HM
    CLASS CORE ;
    FOREIGN DFQRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        ANTENNAGATEAREA 0.126  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.260  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.000 2.300 1.200 ;
        LAYER ME2 ;
        RECT  2.100 0.750 2.300 1.300 ;
        LAYER ME1 ;
        RECT  1.900 0.940 2.340 1.290 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.078  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 3.640 0.840 3.960 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 2.720 1.700 4.370 ;
        RECT  1.300 3.640 1.700 3.960 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.295  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 3.580 3.960 3.960 ;
        RECT  2.320 3.580 3.960 3.780 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 3.960 4.880 4.360 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  2.950 3.080 3.300 3.280 ;
        RECT  2.950 2.260 3.110 3.280 ;
        RECT  2.020 2.260 2.220 2.960 ;
        RECT  1.480 1.780 1.680 2.540 ;
        RECT  0.980 2.260 1.180 3.340 ;
        RECT  0.160 1.520 0.320 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  4.340 -0.140 4.620 0.320 ;
        RECT  3.820 -0.140 4.100 0.320 ;
        RECT  1.100 -0.140 1.380 0.540 ;
        RECT  0.140 -0.140 0.340 0.740 ;
        RECT  0.000 4.660 7.200 4.940 ;
        RECT  3.900 4.480 4.180 4.940 ;
        RECT  1.980 4.300 2.260 4.940 ;
        RECT  0.980 4.240 1.180 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.280 2.700 0.560 3.300 ;
        RECT  0.140 3.100 0.700 3.300 ;
        RECT  0.140 3.100 0.340 4.450 ;
        RECT  0.140 4.250 0.700 4.450 ;
        RECT  2.940 1.480 4.140 1.680 ;
        RECT  2.940 1.480 3.140 1.780 ;
        RECT  3.500 3.080 4.280 3.240 ;
        RECT  2.540 2.720 2.740 3.360 ;
        RECT  1.860 3.180 2.740 3.360 ;
        RECT  4.120 3.460 4.440 3.740 ;
        RECT  1.860 3.180 2.020 4.140 ;
        RECT  1.860 3.980 3.270 4.140 ;
        RECT  3.060 3.980 3.270 4.320 ;
        RECT  4.120 3.080 4.280 4.320 ;
        RECT  3.060 4.160 4.280 4.320 ;
        RECT  1.940 0.620 2.660 0.780 ;
        RECT  2.500 0.800 4.780 0.960 ;
        RECT  4.620 0.800 4.780 1.260 ;
        RECT  2.500 0.620 2.660 1.730 ;
        RECT  2.280 1.530 2.660 1.730 ;
        RECT  1.540 0.300 3.050 0.460 ;
        RECT  2.890 0.300 3.050 0.640 ;
        RECT  2.890 0.480 5.100 0.640 ;
        RECT  0.660 0.460 0.860 0.860 ;
        RECT  1.540 0.300 1.700 0.860 ;
        RECT  0.660 0.700 1.700 0.860 ;
        RECT  4.940 0.480 5.100 1.180 ;
        RECT  4.940 0.970 5.880 1.180 ;
        RECT  0.800 0.700 1.000 1.780 ;
        RECT  0.280 1.060 0.640 1.260 ;
        RECT  1.160 1.460 2.000 1.620 ;
        RECT  0.480 1.060 0.640 2.100 ;
        RECT  1.840 1.460 2.000 2.100 ;
        RECT  1.160 1.460 1.320 2.100 ;
        RECT  0.480 1.940 1.320 2.100 ;
        RECT  1.840 1.940 6.160 2.100 ;
        RECT  5.420 0.340 6.200 0.540 ;
        RECT  2.950 1.140 4.460 1.300 ;
        RECT  4.300 1.140 4.460 1.690 ;
        RECT  6.040 0.340 6.200 1.690 ;
        RECT  4.300 1.530 6.200 1.690 ;
        RECT  4.620 3.080 4.820 3.400 ;
        RECT  6.100 3.120 6.300 3.400 ;
        RECT  4.620 3.240 6.300 3.400 ;
        RECT  5.040 3.240 5.240 4.500 ;
        RECT  6.380 0.310 6.580 1.750 ;
        RECT  3.360 2.700 6.900 2.860 ;
        RECT  3.360 2.700 3.640 2.920 ;
        RECT  6.700 2.700 6.900 4.460 ;
        RECT  5.600 4.260 6.900 4.460 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 3.660 ;
        RECT  5.700 1.140 6.610 3.750 ;
        LAYER VTNH ;
        RECT  0.000 3.660 5.700 4.800 ;
        RECT  6.610 3.660 7.200 4.800 ;
        RECT  0.000 3.750 7.200 4.800 ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END DFQRSM4HM

MACRO DFQRSM2HM
    CLASS CORE ;
    FOREIGN DFQRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.623  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.500 0.970 8.700 1.170 ;
        LAYER ME2 ;
        RECT  8.450 0.800 8.750 1.300 ;
        LAYER ME1 ;
        RECT  8.430 0.940 8.830 1.230 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.430 1.160 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.160 2.560 1.360 ;
        RECT  2.040 1.160 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.510 0.430 11.900 2.100 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.170 0.900 10.890 1.160 ;
        RECT  10.170 0.720 10.330 1.160 ;
        RECT  8.990 0.720 10.330 0.880 ;
        RECT  8.990 0.300 9.150 0.880 ;
        RECT  6.200 0.300 9.150 0.460 ;
        RECT  4.440 1.120 6.360 1.280 ;
        RECT  6.200 0.300 6.360 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  10.990 1.780 11.190 2.540 ;
        RECT  9.910 1.800 10.110 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.880 2.080 6.160 2.540 ;
        RECT  4.440 2.080 4.720 2.540 ;
        RECT  1.560 2.080 1.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  10.830 -0.140 11.030 0.380 ;
        RECT  9.310 -0.140 9.510 0.560 ;
        RECT  4.280 -0.140 4.560 0.320 ;
        RECT  1.700 -0.140 1.980 0.540 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.080 1.520 3.960 1.740 ;
        RECT  2.580 0.620 2.860 0.960 ;
        RECT  2.580 0.800 5.280 0.960 ;
        RECT  2.720 0.800 2.900 1.740 ;
        RECT  2.460 1.540 2.900 1.740 ;
        RECT  2.140 0.300 3.280 0.460 ;
        RECT  3.120 0.300 3.280 0.640 ;
        RECT  3.120 0.480 6.040 0.640 ;
        RECT  1.260 0.340 1.460 0.860 ;
        RECT  2.140 0.300 2.300 0.860 ;
        RECT  1.260 0.700 2.300 0.860 ;
        RECT  5.760 0.480 6.040 0.960 ;
        RECT  1.400 0.700 1.600 1.600 ;
        RECT  1.220 1.440 1.600 1.600 ;
        RECT  0.140 0.340 0.340 0.640 ;
        RECT  0.140 0.480 0.980 0.640 ;
        RECT  0.100 1.550 0.980 1.750 ;
        RECT  0.820 0.480 0.980 1.920 ;
        RECT  0.820 1.760 2.250 1.920 ;
        RECT  4.120 1.760 5.040 1.920 ;
        RECT  5.560 1.760 7.010 1.920 ;
        RECT  2.090 1.760 2.250 2.100 ;
        RECT  4.880 1.760 5.040 2.100 ;
        RECT  4.120 1.760 4.280 2.100 ;
        RECT  2.090 1.940 4.280 2.100 ;
        RECT  5.560 1.760 5.720 2.100 ;
        RECT  4.880 1.940 5.720 2.100 ;
        RECT  3.300 1.120 4.280 1.320 ;
        RECT  4.120 1.120 4.280 1.600 ;
        RECT  6.520 0.620 6.800 1.600 ;
        RECT  4.120 1.440 7.330 1.600 ;
        RECT  5.200 1.440 5.400 1.780 ;
        RECT  7.170 1.440 7.330 1.800 ;
        RECT  7.630 0.620 8.610 0.780 ;
        RECT  8.110 0.620 8.270 1.720 ;
        RECT  8.110 1.440 9.690 1.600 ;
        RECT  8.110 1.440 8.480 1.720 ;
        RECT  7.040 0.620 7.320 1.250 ;
        RECT  7.040 1.050 7.850 1.250 ;
        RECT  8.640 1.760 9.730 1.920 ;
        RECT  7.690 1.050 7.850 2.100 ;
        RECT  8.640 1.760 8.800 2.100 ;
        RECT  7.690 1.940 8.800 2.100 ;
        RECT  9.450 1.760 9.730 2.100 ;
        RECT  9.850 0.320 10.650 0.520 ;
        RECT  10.490 0.320 10.650 0.740 ;
        RECT  10.490 0.580 11.310 0.740 ;
        RECT  8.990 1.040 10.010 1.240 ;
        RECT  9.850 1.040 10.010 1.620 ;
        RECT  11.150 0.580 11.310 1.620 ;
        RECT  9.850 1.420 11.310 1.620 ;
        RECT  10.470 1.420 10.670 1.970 ;
        LAYER VTPH ;
        RECT  0.550 1.080 1.750 2.400 ;
        RECT  8.910 1.070 9.850 2.400 ;
        RECT  0.000 1.140 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.070 ;
        RECT  0.000 0.000 8.910 1.080 ;
        RECT  0.000 0.000 0.550 1.140 ;
        RECT  1.750 0.000 8.910 1.140 ;
        RECT  9.850 0.000 12.000 1.140 ;
    END
END DFQRSM2HM

MACRO DFQRSM1HM
    CLASS CORE ;
    FOREIGN DFQRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.124  LAYER ME1  ;
        ANTENNAGATEAREA 0.124  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.903  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.500 0.970 8.700 1.170 ;
        LAYER ME2 ;
        RECT  8.450 0.800 8.750 1.300 ;
        LAYER ME1 ;
        RECT  8.430 0.940 8.830 1.230 ;
        END
    END SB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.430 1.160 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.103  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.160 2.560 1.360 ;
        RECT  2.040 1.160 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.313  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.530 0.360 11.900 1.970 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.170 0.900 10.890 1.160 ;
        RECT  10.170 0.720 10.330 1.160 ;
        RECT  8.990 0.720 10.330 0.880 ;
        RECT  8.990 0.300 9.150 0.880 ;
        RECT  6.200 0.300 9.150 0.460 ;
        RECT  4.440 1.120 6.360 1.280 ;
        RECT  6.200 0.300 6.360 1.280 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.000 2.540 ;
        RECT  10.990 1.780 11.190 2.540 ;
        RECT  9.910 1.800 10.110 2.540 ;
        RECT  8.960 2.080 9.240 2.540 ;
        RECT  5.880 2.080 6.160 2.540 ;
        RECT  4.440 2.080 4.720 2.540 ;
        RECT  1.560 2.080 1.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.000 0.140 ;
        RECT  10.830 -0.140 11.030 0.380 ;
        RECT  9.310 -0.140 9.510 0.560 ;
        RECT  4.280 -0.140 4.560 0.320 ;
        RECT  1.700 -0.140 1.980 0.540 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.080 1.520 3.960 1.740 ;
        RECT  2.580 0.620 2.860 0.960 ;
        RECT  2.580 0.800 5.280 0.960 ;
        RECT  2.720 0.800 2.900 1.740 ;
        RECT  2.460 1.540 2.900 1.740 ;
        RECT  2.140 0.300 3.280 0.460 ;
        RECT  3.120 0.300 3.280 0.640 ;
        RECT  3.120 0.480 6.040 0.640 ;
        RECT  1.260 0.340 1.460 0.860 ;
        RECT  2.140 0.300 2.300 0.860 ;
        RECT  1.260 0.700 2.300 0.860 ;
        RECT  5.760 0.480 6.040 0.960 ;
        RECT  1.400 0.700 1.600 1.600 ;
        RECT  1.220 1.440 1.600 1.600 ;
        RECT  0.140 0.340 0.340 0.640 ;
        RECT  0.140 0.480 0.980 0.640 ;
        RECT  0.100 1.550 0.980 1.750 ;
        RECT  0.820 0.480 0.980 1.920 ;
        RECT  0.820 1.760 2.250 1.920 ;
        RECT  4.120 1.760 5.040 1.920 ;
        RECT  5.560 1.760 6.950 1.920 ;
        RECT  2.090 1.760 2.250 2.100 ;
        RECT  4.880 1.760 5.040 2.100 ;
        RECT  4.120 1.760 4.280 2.100 ;
        RECT  2.090 1.940 4.280 2.100 ;
        RECT  5.560 1.760 5.720 2.100 ;
        RECT  4.880 1.940 5.720 2.100 ;
        RECT  3.300 1.120 4.280 1.320 ;
        RECT  4.120 1.120 4.280 1.600 ;
        RECT  6.520 0.620 6.800 1.600 ;
        RECT  4.120 1.440 7.350 1.600 ;
        RECT  7.150 1.440 7.350 1.720 ;
        RECT  5.200 1.440 5.400 1.780 ;
        RECT  7.630 0.620 8.610 0.780 ;
        RECT  8.110 0.620 8.270 1.720 ;
        RECT  8.110 1.440 9.690 1.600 ;
        RECT  8.110 1.440 8.480 1.720 ;
        RECT  7.040 0.620 7.320 1.250 ;
        RECT  7.040 1.050 7.850 1.250 ;
        RECT  8.640 1.760 9.730 1.920 ;
        RECT  7.690 1.050 7.850 2.100 ;
        RECT  8.640 1.760 8.800 2.100 ;
        RECT  7.690 1.940 8.800 2.100 ;
        RECT  9.450 1.760 9.730 2.100 ;
        RECT  9.850 0.320 10.650 0.520 ;
        RECT  10.490 0.320 10.650 0.740 ;
        RECT  10.490 0.580 11.310 0.740 ;
        RECT  8.990 1.040 10.010 1.240 ;
        RECT  9.850 1.040 10.010 1.620 ;
        RECT  11.150 0.580 11.310 1.620 ;
        RECT  9.850 1.420 11.310 1.620 ;
        RECT  10.470 1.420 10.670 2.080 ;
        LAYER VTPH ;
        RECT  0.550 1.080 1.750 2.400 ;
        RECT  8.910 1.070 9.850 2.400 ;
        RECT  0.000 1.140 12.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.000 1.070 ;
        RECT  0.000 0.000 8.910 1.080 ;
        RECT  0.000 0.000 0.550 1.140 ;
        RECT  1.750 0.000 8.910 1.140 ;
        RECT  9.850 0.000 12.000 1.140 ;
    END
END DFQRSM1HM

MACRO DFQRM8HM
    CLASS CORE ;
    FOREIGN DFQRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.254  LAYER ME1  ;
        ANTENNAGATEAREA 0.254  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.709  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.700 1.800 7.900 2.000 ;
        LAYER ME2 ;
        RECT  7.600 1.640 8.000 2.000 ;
        LAYER ME1 ;
        RECT  7.490 1.760 8.130 2.100 ;
        RECT  6.560 1.760 8.130 1.920 ;
        RECT  5.380 1.940 6.720 2.100 ;
        RECT  6.560 1.760 6.720 2.100 ;
        RECT  5.380 1.540 5.540 2.100 ;
        RECT  4.620 1.540 5.540 1.700 ;
        RECT  4.620 1.540 4.780 2.020 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        ANTENNAGATEAREA 0.120  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.250  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.380 1.090 2.580 1.290 ;
        LAYER ME2 ;
        RECT  2.360 1.000 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.300 1.000 2.650 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.420 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.760 0.380 11.960 2.100 ;
        RECT  10.720 0.900 11.960 1.100 ;
        RECT  10.720 0.380 10.920 2.080 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  12.280 1.480 12.480 2.540 ;
        RECT  11.240 1.480 11.440 2.540 ;
        RECT  10.200 1.480 10.400 2.540 ;
        RECT  9.840 1.480 10.040 2.540 ;
        RECT  8.710 1.760 8.910 2.540 ;
        RECT  8.290 1.760 8.490 2.540 ;
        RECT  6.960 2.080 7.240 2.540 ;
        RECT  4.940 1.860 5.220 2.540 ;
        RECT  3.700 1.860 3.980 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  12.280 -0.140 12.480 0.660 ;
        RECT  11.240 -0.140 11.440 0.660 ;
        RECT  10.180 -0.140 10.340 0.420 ;
        RECT  8.290 -0.140 8.450 0.420 ;
        RECT  6.700 -0.140 6.980 0.320 ;
        RECT  4.020 -0.140 4.300 0.320 ;
        RECT  1.660 -0.140 1.860 0.380 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.440 0.340 0.860 ;
        RECT  0.140 0.700 0.840 0.860 ;
        RECT  0.680 1.000 1.180 1.200 ;
        RECT  0.680 0.700 0.840 1.920 ;
        RECT  0.100 1.720 0.840 1.920 ;
        RECT  0.100 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  1.100 1.940 3.200 2.100 ;
        RECT  3.140 1.500 4.420 1.660 ;
        RECT  3.140 1.500 3.340 1.780 ;
        RECT  4.220 1.500 4.420 1.780 ;
        RECT  2.540 0.620 2.980 0.840 ;
        RECT  2.810 0.800 4.600 0.960 ;
        RECT  2.810 0.620 2.970 1.780 ;
        RECT  2.460 1.620 2.970 1.780 ;
        RECT  5.080 0.620 5.360 1.340 ;
        RECT  3.180 1.180 5.860 1.340 ;
        RECT  5.700 1.180 5.860 1.760 ;
        RECT  2.210 0.300 3.800 0.460 ;
        RECT  4.540 0.300 5.680 0.460 ;
        RECT  3.640 0.300 3.800 0.640 ;
        RECT  1.180 0.340 1.380 0.700 ;
        RECT  4.540 0.300 4.700 0.640 ;
        RECT  3.640 0.480 4.700 0.640 ;
        RECT  2.210 0.300 2.380 0.700 ;
        RECT  1.180 0.540 2.380 0.700 ;
        RECT  5.520 0.300 5.680 1.020 ;
        RECT  5.520 0.840 6.590 1.020 ;
        RECT  6.390 0.840 6.590 1.280 ;
        RECT  1.900 0.540 2.060 1.600 ;
        RECT  1.040 1.440 2.060 1.600 ;
        RECT  5.840 0.300 6.040 0.680 ;
        RECT  5.840 0.520 7.550 0.680 ;
        RECT  7.390 0.520 7.550 1.200 ;
        RECT  7.390 1.000 8.910 1.200 ;
        RECT  6.750 0.520 6.910 1.600 ;
        RECT  6.200 1.440 6.910 1.600 ;
        RECT  6.200 1.440 6.400 1.720 ;
        RECT  8.710 0.300 9.990 0.460 ;
        RECT  7.730 0.320 7.890 0.780 ;
        RECT  8.710 0.300 8.910 0.780 ;
        RECT  7.730 0.610 8.910 0.780 ;
        RECT  9.790 0.300 9.990 0.840 ;
        RECT  9.230 1.080 10.510 1.280 ;
        RECT  7.070 0.960 7.230 1.600 ;
        RECT  7.070 1.440 9.510 1.600 ;
        RECT  9.230 0.620 9.510 1.930 ;
        LAYER VTPH ;
        RECT  5.720 1.080 8.520 2.400 ;
        RECT  0.520 1.080 2.170 2.400 ;
        RECT  0.000 1.140 2.170 2.400 ;
        RECT  3.190 1.140 12.800 2.400 ;
        RECT  0.000 1.170 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.080 ;
        RECT  0.000 0.000 0.520 1.140 ;
        RECT  2.170 0.000 5.720 1.140 ;
        RECT  8.520 0.000 12.800 1.140 ;
        RECT  2.170 0.000 3.190 1.170 ;
    END
END DFQRM8HM

MACRO DFQRM4HM
    CLASS CORE ;
    FOREIGN DFQRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.254  LAYER ME1  ;
        ANTENNAGATEAREA 0.254  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.627  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.650 1.800 7.850 2.000 ;
        LAYER ME2 ;
        RECT  7.550 1.640 7.950 2.000 ;
        LAYER ME1 ;
        RECT  7.460 1.760 8.100 2.100 ;
        RECT  6.600 1.760 8.100 1.920 ;
        RECT  5.350 1.900 6.760 2.100 ;
        RECT  5.350 1.540 5.510 2.100 ;
        RECT  4.590 1.540 5.510 1.700 ;
        RECT  4.590 1.540 4.750 2.020 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.420 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.160 2.480 1.360 ;
        RECT  2.100 1.160 2.300 1.560 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.690 0.420 10.890 2.100 ;
        RECT  10.500 1.200 10.890 1.650 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.210 1.480 11.410 2.540 ;
        RECT  10.120 1.460 10.320 2.540 ;
        RECT  9.760 1.590 9.960 2.540 ;
        RECT  8.680 1.760 8.880 2.540 ;
        RECT  8.260 1.760 8.460 2.540 ;
        RECT  6.930 2.080 7.210 2.540 ;
        RECT  4.910 1.860 5.190 2.540 ;
        RECT  3.660 1.860 3.960 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.210 -0.140 11.410 0.660 ;
        RECT  10.150 -0.140 10.310 0.420 ;
        RECT  8.160 -0.140 8.440 0.500 ;
        RECT  7.100 -0.140 7.380 0.500 ;
        RECT  3.980 -0.140 4.260 0.320 ;
        RECT  1.660 -0.140 1.860 0.560 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 0.340 0.860 ;
        RECT  0.140 0.660 0.840 0.860 ;
        RECT  0.680 1.040 1.240 1.240 ;
        RECT  0.680 0.660 0.840 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  0.140 1.760 0.340 2.100 ;
        RECT  1.100 1.940 3.160 2.100 ;
        RECT  3.060 1.500 4.430 1.680 ;
        RECT  4.150 1.500 4.430 1.700 ;
        RECT  3.060 1.500 3.340 1.720 ;
        RECT  2.460 0.620 2.820 0.780 ;
        RECT  2.640 0.800 4.560 0.960 ;
        RECT  2.640 0.620 2.820 1.780 ;
        RECT  2.460 1.580 2.820 1.780 ;
        RECT  5.050 0.620 5.330 1.340 ;
        RECT  3.140 1.180 5.870 1.340 ;
        RECT  5.670 1.180 5.870 1.720 ;
        RECT  2.020 0.300 3.760 0.460 ;
        RECT  4.420 0.300 5.650 0.460 ;
        RECT  3.600 0.300 3.760 0.640 ;
        RECT  4.420 0.300 4.580 0.640 ;
        RECT  3.600 0.480 4.580 0.640 ;
        RECT  1.180 0.300 1.380 0.880 ;
        RECT  5.490 0.300 5.650 1.020 ;
        RECT  2.020 0.300 2.190 0.880 ;
        RECT  1.180 0.720 2.190 0.880 ;
        RECT  5.490 0.840 6.560 1.020 ;
        RECT  6.360 0.840 6.560 1.280 ;
        RECT  1.590 0.720 1.790 1.600 ;
        RECT  1.100 1.440 1.790 1.600 ;
        RECT  5.810 0.300 6.010 0.680 ;
        RECT  5.810 0.520 6.880 0.680 ;
        RECT  6.720 0.660 7.560 0.820 ;
        RECT  7.400 0.660 7.560 1.200 ;
        RECT  7.400 1.000 8.580 1.200 ;
        RECT  6.720 0.520 6.880 1.600 ;
        RECT  6.170 1.440 6.880 1.600 ;
        RECT  6.170 1.440 6.370 1.720 ;
        RECT  8.680 0.300 9.960 0.460 ;
        RECT  7.640 0.320 7.920 0.520 ;
        RECT  7.760 0.320 7.920 0.820 ;
        RECT  8.680 0.300 8.880 0.820 ;
        RECT  7.760 0.660 8.880 0.820 ;
        RECT  9.760 0.300 9.960 0.840 ;
        RECT  9.200 0.620 9.480 1.280 ;
        RECT  9.200 1.080 10.230 1.280 ;
        RECT  7.040 0.980 7.240 1.600 ;
        RECT  9.200 0.620 9.440 1.600 ;
        RECT  7.040 1.440 9.440 1.600 ;
        RECT  9.240 0.620 9.440 1.880 ;
        LAYER VTPH ;
        RECT  5.720 1.080 8.900 2.400 ;
        RECT  0.430 1.080 2.170 2.400 ;
        RECT  0.000 1.140 2.170 2.400 ;
        RECT  3.270 1.140 11.600 2.400 ;
        RECT  0.000 1.170 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.080 ;
        RECT  0.000 0.000 0.430 1.140 ;
        RECT  2.170 0.000 5.720 1.140 ;
        RECT  8.900 0.000 11.600 1.140 ;
        RECT  2.170 0.000 3.270 1.170 ;
    END
END DFQRM4HM

MACRO DFQRM2HM
    CLASS CORE ;
    FOREIGN DFQRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.146  LAYER ME1  ;
        ANTENNAGATEAREA 0.146  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 15.522  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.520 1.800 7.720 2.000 ;
        LAYER ME2 ;
        RECT  7.300 1.640 7.820 2.000 ;
        LAYER ME1 ;
        RECT  7.460 1.760 7.780 2.100 ;
        RECT  6.600 1.760 7.780 1.920 ;
        RECT  5.370 1.900 6.760 2.100 ;
        RECT  5.370 1.540 5.530 2.100 ;
        RECT  4.610 1.540 5.530 1.700 ;
        RECT  4.610 1.540 4.770 2.020 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.420 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.160 2.530 1.360 ;
        RECT  2.100 1.160 2.300 1.570 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.260 0.380 9.500 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.740 1.440 8.940 2.540 ;
        RECT  6.950 2.080 7.230 2.540 ;
        RECT  4.930 1.860 5.210 2.540 ;
        RECT  3.680 1.860 3.980 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.740 -0.140 8.940 0.700 ;
        RECT  7.070 -0.140 7.350 0.500 ;
        RECT  4.000 -0.140 4.280 0.320 ;
        RECT  1.660 -0.140 1.860 0.560 ;
        RECT  0.660 -0.140 0.860 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 0.340 0.900 ;
        RECT  0.140 0.720 0.840 0.900 ;
        RECT  0.680 1.040 1.240 1.240 ;
        RECT  0.680 0.720 0.840 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  0.140 1.760 0.340 2.100 ;
        RECT  1.100 1.940 3.180 2.100 ;
        RECT  3.080 1.500 4.450 1.680 ;
        RECT  4.170 1.500 4.450 1.700 ;
        RECT  3.080 1.500 3.360 1.720 ;
        RECT  2.540 0.620 2.860 0.840 ;
        RECT  2.690 0.800 4.700 0.960 ;
        RECT  2.690 0.620 2.850 1.780 ;
        RECT  2.480 1.580 2.850 1.780 ;
        RECT  5.070 0.620 5.350 1.340 ;
        RECT  3.160 1.180 5.890 1.340 ;
        RECT  5.690 1.180 5.890 1.720 ;
        RECT  2.020 0.300 3.460 0.460 ;
        RECT  4.440 0.300 5.670 0.460 ;
        RECT  3.300 0.300 3.460 0.640 ;
        RECT  4.440 0.300 4.600 0.640 ;
        RECT  3.300 0.480 4.600 0.640 ;
        RECT  1.180 0.300 1.380 0.880 ;
        RECT  5.510 0.300 5.670 1.020 ;
        RECT  2.020 0.300 2.190 0.880 ;
        RECT  1.180 0.720 2.190 0.880 ;
        RECT  5.510 0.840 6.580 1.020 ;
        RECT  6.380 0.840 6.580 1.280 ;
        RECT  1.590 0.720 1.790 1.600 ;
        RECT  1.040 1.440 1.790 1.600 ;
        RECT  5.830 0.300 6.030 0.680 ;
        RECT  5.830 0.520 6.900 0.680 ;
        RECT  6.740 0.660 8.040 0.820 ;
        RECT  7.840 0.660 8.040 1.240 ;
        RECT  6.740 0.520 6.900 1.600 ;
        RECT  6.190 1.440 6.900 1.600 ;
        RECT  6.190 1.440 6.390 1.720 ;
        RECT  7.940 0.340 8.360 0.500 ;
        RECT  8.200 1.000 9.080 1.200 ;
        RECT  7.060 0.980 7.260 1.600 ;
        RECT  7.060 1.440 8.360 1.600 ;
        RECT  8.200 0.340 8.360 2.000 ;
        LAYER VTPH ;
        RECT  5.580 1.080 8.300 2.400 ;
        RECT  0.430 1.080 2.170 2.400 ;
        RECT  0.000 1.140 2.170 2.400 ;
        RECT  3.170 1.140 9.600 2.400 ;
        RECT  0.000 1.170 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.080 ;
        RECT  0.000 0.000 0.430 1.140 ;
        RECT  2.170 0.000 5.580 1.140 ;
        RECT  8.300 0.000 9.600 1.140 ;
        RECT  2.170 0.000 3.170 1.170 ;
    END
END DFQRM2HM

MACRO DFQRM1HM
    CLASS CORE ;
    FOREIGN DFQRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.210  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.200 1.090 2.400 1.290 ;
        LAYER ME2 ;
        RECT  2.100 1.000 2.400 1.560 ;
        LAYER ME1 ;
        RECT  2.150 1.010 2.440 1.400 ;
        END
    END D
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        ANTENNAGATEAREA 0.119  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 19.172  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  7.530 1.760 7.730 1.960 ;
        LAYER ME2 ;
        RECT  7.470 1.640 7.900 2.000 ;
        LAYER ME1 ;
        RECT  7.470 1.760 7.810 2.100 ;
        RECT  6.250 1.760 7.810 1.920 ;
        RECT  5.390 1.900 6.410 2.100 ;
        RECT  5.390 1.540 5.550 2.100 ;
        RECT  4.630 1.540 5.550 1.700 ;
        RECT  4.630 1.540 4.790 2.020 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.100 0.420 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.150 1.840 9.500 2.040 ;
        RECT  9.300 0.420 9.500 2.040 ;
        RECT  9.150 0.420 9.500 0.620 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.670 1.800 8.870 2.540 ;
        RECT  7.030 2.080 7.310 2.540 ;
        RECT  4.950 1.860 5.230 2.540 ;
        RECT  3.700 1.860 4.000 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.660 -0.140 8.870 0.630 ;
        RECT  7.050 -0.140 7.330 0.500 ;
        RECT  4.020 -0.140 4.300 0.320 ;
        RECT  1.660 -0.140 1.860 0.380 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 0.340 0.840 ;
        RECT  0.140 0.660 0.840 0.840 ;
        RECT  0.680 1.000 1.240 1.200 ;
        RECT  0.680 0.660 0.840 1.920 ;
        RECT  0.140 1.760 1.260 1.920 ;
        RECT  1.100 1.760 1.260 2.100 ;
        RECT  0.140 1.760 0.340 2.100 ;
        RECT  1.100 1.940 3.200 2.100 ;
        RECT  3.100 1.500 4.470 1.680 ;
        RECT  4.190 1.500 4.470 1.700 ;
        RECT  3.100 1.500 3.380 1.720 ;
        RECT  2.540 0.620 2.820 0.840 ;
        RECT  2.640 0.800 4.720 0.960 ;
        RECT  2.640 0.620 2.820 1.780 ;
        RECT  2.460 1.620 2.820 1.780 ;
        RECT  5.090 0.620 5.370 1.340 ;
        RECT  3.180 1.180 5.910 1.340 ;
        RECT  5.710 1.180 5.910 1.720 ;
        RECT  2.210 0.300 3.800 0.460 ;
        RECT  4.460 0.300 5.690 0.460 ;
        RECT  3.640 0.300 3.800 0.640 ;
        RECT  1.180 0.300 1.380 0.700 ;
        RECT  4.460 0.300 4.620 0.640 ;
        RECT  3.640 0.480 4.620 0.640 ;
        RECT  2.210 0.300 2.380 0.700 ;
        RECT  1.180 0.540 2.380 0.700 ;
        RECT  5.530 0.300 5.690 1.020 ;
        RECT  5.530 0.860 6.570 1.020 ;
        RECT  6.370 0.860 6.570 1.280 ;
        RECT  1.750 0.540 1.950 1.600 ;
        RECT  1.100 1.440 1.950 1.600 ;
        RECT  5.850 0.300 6.050 0.680 ;
        RECT  5.850 0.520 6.890 0.680 ;
        RECT  6.730 0.660 8.030 0.820 ;
        RECT  7.830 0.660 8.030 1.180 ;
        RECT  6.730 0.520 6.890 1.600 ;
        RECT  6.170 1.440 6.890 1.600 ;
        RECT  7.930 0.340 8.410 0.500 ;
        RECT  8.250 1.080 9.090 1.280 ;
        RECT  7.050 1.000 7.250 1.600 ;
        RECT  7.050 1.440 8.410 1.600 ;
        RECT  8.250 0.340 8.410 2.100 ;
        RECT  8.170 1.440 8.410 2.100 ;
        LAYER VTPH ;
        RECT  5.600 1.080 8.140 2.400 ;
        RECT  0.430 1.080 1.640 2.400 ;
        RECT  0.000 1.140 1.640 2.400 ;
        RECT  3.190 1.140 9.600 2.400 ;
        RECT  0.000 1.170 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.080 ;
        RECT  0.000 0.000 0.430 1.140 ;
        RECT  1.640 0.000 5.600 1.140 ;
        RECT  8.140 0.000 9.600 1.140 ;
        RECT  1.640 0.000 3.190 1.170 ;
    END
END DFQRM1HM

MACRO DFQM8HM
    CLASS CORE ;
    FOREIGN DFQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        ANTENNAGATEAREA 0.131  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.783  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.460 1.040 2.660 1.240 ;
        LAYER ME2 ;
        RECT  2.460 0.750 2.700 1.300 ;
        LAYER ME1 ;
        RECT  2.420 0.940 2.660 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 0.430 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.339  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.020 1.460 9.220 2.100 ;
        RECT  6.940 0.770 9.220 0.940 ;
        RECT  9.020 0.430 9.220 0.940 ;
        RECT  6.940 1.460 9.220 1.660 ;
        RECT  8.500 0.770 8.700 1.660 ;
        RECT  7.980 1.460 8.200 2.100 ;
        RECT  7.980 0.430 8.180 0.940 ;
        RECT  6.940 1.460 7.140 2.100 ;
        RECT  6.940 0.430 7.140 0.940 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.500 1.840 8.700 2.540 ;
        RECT  7.460 1.840 7.660 2.540 ;
        RECT  5.900 1.470 6.100 2.540 ;
        RECT  3.480 2.020 3.680 2.540 ;
        RECT  1.560 2.080 1.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.500 -0.140 8.700 0.560 ;
        RECT  7.460 -0.140 7.660 0.560 ;
        RECT  5.900 -0.140 6.100 0.380 ;
        RECT  3.480 -0.140 3.760 0.320 ;
        RECT  1.740 -0.140 1.940 0.640 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.560 0.620 2.980 0.780 ;
        RECT  3.820 1.120 4.020 1.540 ;
        RECT  2.820 1.380 4.020 1.540 ;
        RECT  2.820 0.620 2.980 1.720 ;
        RECT  2.400 1.560 2.980 1.720 ;
        RECT  3.340 0.800 4.440 0.960 ;
        RECT  3.340 0.800 3.540 1.220 ;
        RECT  4.240 0.620 4.440 1.780 ;
        RECT  4.180 0.800 4.440 1.780 ;
        RECT  0.140 0.440 0.340 0.860 ;
        RECT  0.140 0.700 1.020 0.860 ;
        RECT  0.860 0.700 1.020 1.920 ;
        RECT  0.100 1.720 1.020 1.920 ;
        RECT  3.140 1.700 4.000 1.860 ;
        RECT  0.100 1.760 2.160 1.920 ;
        RECT  2.000 1.760 2.160 2.100 ;
        RECT  3.840 1.700 4.000 2.100 ;
        RECT  3.140 1.700 3.300 2.100 ;
        RECT  2.000 1.940 3.300 2.100 ;
        RECT  3.840 1.940 4.560 2.100 ;
        RECT  2.100 0.300 3.300 0.460 ;
        RECT  3.920 0.300 5.380 0.460 ;
        RECT  3.140 0.300 3.300 0.640 ;
        RECT  3.920 0.300 4.080 0.640 ;
        RECT  3.140 0.480 4.080 0.640 ;
        RECT  1.220 0.450 1.580 0.650 ;
        RECT  2.100 0.300 2.260 0.960 ;
        RECT  1.420 0.800 2.260 0.960 ;
        RECT  1.420 0.450 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  5.180 0.300 5.380 1.720 ;
        RECT  5.540 1.110 6.240 1.310 ;
        RECT  4.720 0.620 4.920 2.100 ;
        RECT  5.540 1.110 5.700 2.100 ;
        RECT  4.720 1.940 5.700 2.100 ;
        RECT  5.540 0.680 6.660 0.880 ;
        RECT  6.460 1.100 8.240 1.300 ;
        RECT  6.460 0.430 6.660 2.090 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.720 2.400 ;
        RECT  0.000 1.140 2.950 2.400 ;
        RECT  5.160 1.140 9.600 2.400 ;
        RECT  0.000 1.200 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.720 0.000 9.600 1.140 ;
        RECT  2.950 0.000 5.160 1.200 ;
    END
END DFQM8HM

MACRO DFQM4HM
    CLASS CORE ;
    FOREIGN DFQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.655  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.460 1.040 2.660 1.240 ;
        LAYER ME2 ;
        RECT  2.460 0.750 2.700 1.300 ;
        LAYER ME1 ;
        RECT  2.420 0.940 2.660 1.400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 0.430 1.560 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.843  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.010 1.460 8.300 2.100 ;
        RECT  8.030 0.430 8.300 2.100 ;
        RECT  6.970 0.770 8.300 0.940 ;
        RECT  8.010 0.430 8.300 0.940 ;
        RECT  6.970 1.460 8.300 1.660 ;
        RECT  6.970 1.460 7.170 2.100 ;
        RECT  6.970 0.430 7.170 0.940 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.490 1.840 7.690 2.540 ;
        RECT  5.930 1.470 6.130 2.540 ;
        RECT  3.480 2.020 3.680 2.540 ;
        RECT  1.560 2.080 1.840 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.490 -0.140 7.690 0.560 ;
        RECT  5.930 -0.140 6.130 0.380 ;
        RECT  3.480 -0.140 3.760 0.320 ;
        RECT  1.740 -0.140 1.940 0.640 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.560 0.620 2.980 0.780 ;
        RECT  3.820 1.120 4.020 1.540 ;
        RECT  2.820 1.380 4.020 1.540 ;
        RECT  2.820 0.620 2.980 1.720 ;
        RECT  2.430 1.560 2.980 1.720 ;
        RECT  3.340 0.800 4.440 0.960 ;
        RECT  3.340 0.800 3.540 1.220 ;
        RECT  4.240 0.620 4.440 1.780 ;
        RECT  4.180 0.800 4.440 1.780 ;
        RECT  0.140 0.350 0.340 0.860 ;
        RECT  0.140 0.700 1.020 0.860 ;
        RECT  0.860 0.700 1.020 1.920 ;
        RECT  0.100 1.720 1.020 1.920 ;
        RECT  3.140 1.700 4.000 1.860 ;
        RECT  0.100 1.760 2.160 1.920 ;
        RECT  2.000 1.760 2.160 2.100 ;
        RECT  3.840 1.700 4.000 2.100 ;
        RECT  3.140 1.700 3.300 2.100 ;
        RECT  2.000 1.940 3.300 2.100 ;
        RECT  3.840 1.940 4.560 2.100 ;
        RECT  2.100 0.300 3.300 0.460 ;
        RECT  3.920 0.300 5.410 0.460 ;
        RECT  3.140 0.300 3.300 0.640 ;
        RECT  1.220 0.390 1.580 0.590 ;
        RECT  3.920 0.300 4.080 0.640 ;
        RECT  3.140 0.480 4.080 0.640 ;
        RECT  2.100 0.300 2.260 0.960 ;
        RECT  1.420 0.800 2.260 0.960 ;
        RECT  1.420 0.390 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  5.250 0.300 5.410 1.720 ;
        RECT  5.570 1.100 6.280 1.300 ;
        RECT  4.720 0.620 4.950 2.100 ;
        RECT  5.570 1.100 5.730 2.100 ;
        RECT  4.720 1.940 5.730 2.100 ;
        RECT  5.570 0.680 6.690 0.880 ;
        RECT  6.490 1.100 7.690 1.300 ;
        RECT  6.490 0.430 6.690 2.090 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.720 2.400 ;
        RECT  0.000 1.140 2.950 2.400 ;
        RECT  5.200 1.140 8.400 2.400 ;
        RECT  0.000 1.200 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.720 0.000 8.400 1.140 ;
        RECT  2.950 0.000 5.200 1.200 ;
    END
END DFQM4HM

MACRO DFQM2HM
    CLASS CORE ;
    FOREIGN DFQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 0.360 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.240 2.700 1.440 ;
        RECT  2.420 1.120 2.700 1.440 ;
        RECT  2.040 1.240 2.360 1.500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.020 1.460 7.900 1.660 ;
        RECT  7.700 0.760 7.900 1.660 ;
        RECT  7.020 0.760 7.900 0.920 ;
        RECT  7.020 0.430 7.230 0.920 ;
        RECT  7.020 1.460 7.220 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.540 1.840 7.740 2.540 ;
        RECT  6.020 1.680 6.220 2.540 ;
        RECT  3.620 2.080 3.900 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.540 -0.140 7.740 0.600 ;
        RECT  5.930 -0.140 6.130 0.380 ;
        RECT  3.560 -0.140 3.840 0.320 ;
        RECT  1.740 -0.140 1.940 0.600 ;
        RECT  0.620 -0.140 0.900 0.550 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.580 0.620 3.020 0.780 ;
        RECT  2.860 1.440 4.180 1.600 ;
        RECT  3.980 1.120 4.180 1.600 ;
        RECT  2.860 0.620 3.020 1.760 ;
        RECT  2.560 1.600 3.020 1.760 ;
        RECT  4.370 0.620 4.580 0.960 ;
        RECT  3.500 0.800 4.580 0.960 ;
        RECT  3.500 0.800 3.700 1.280 ;
        RECT  4.380 0.620 4.580 1.780 ;
        RECT  0.140 0.350 0.340 0.890 ;
        RECT  0.140 0.730 1.020 0.890 ;
        RECT  0.860 0.730 1.020 1.920 ;
        RECT  0.140 1.750 1.020 1.920 ;
        RECT  0.140 1.760 2.270 1.920 ;
        RECT  3.290 1.760 4.220 1.920 ;
        RECT  2.110 1.760 2.270 2.100 ;
        RECT  4.060 1.760 4.220 2.100 ;
        RECT  0.140 1.750 0.340 2.070 ;
        RECT  3.290 1.760 3.450 2.100 ;
        RECT  2.110 1.940 3.450 2.100 ;
        RECT  4.060 1.940 4.720 2.100 ;
        RECT  2.130 0.300 3.340 0.460 ;
        RECT  4.050 0.300 5.450 0.460 ;
        RECT  3.180 0.300 3.340 0.640 ;
        RECT  1.220 0.340 1.580 0.540 ;
        RECT  4.050 0.300 4.210 0.640 ;
        RECT  3.180 0.480 4.210 0.640 ;
        RECT  2.130 0.300 2.300 0.990 ;
        RECT  1.420 0.830 2.300 0.990 ;
        RECT  5.290 0.300 5.450 1.760 ;
        RECT  1.420 0.340 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  5.290 1.480 5.500 1.760 ;
        RECT  5.670 1.160 6.360 1.360 ;
        RECT  4.890 0.620 5.090 2.100 ;
        RECT  5.670 1.160 5.830 2.100 ;
        RECT  4.890 1.940 5.830 2.100 ;
        RECT  5.660 0.680 6.740 0.880 ;
        RECT  6.540 1.100 7.410 1.300 ;
        RECT  6.540 0.370 6.740 1.850 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.730 2.400 ;
        RECT  0.000 1.140 3.730 2.400 ;
        RECT  5.320 1.140 8.000 2.400 ;
        RECT  0.000 1.200 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.730 0.000 8.000 1.140 ;
        RECT  3.730 0.000 5.320 1.200 ;
    END
END DFQM2HM

MACRO DFQM1HM
    CLASS CORE ;
    FOREIGN DFQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.140 0.360 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.240 2.700 1.440 ;
        RECT  2.420 1.120 2.700 1.440 ;
        RECT  2.040 1.240 2.360 1.500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.020 1.500 7.900 1.680 ;
        RECT  7.700 0.770 7.900 1.680 ;
        RECT  7.020 0.770 7.900 0.940 ;
        RECT  7.020 1.500 7.220 2.100 ;
        RECT  7.020 0.300 7.220 0.940 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.540 1.840 7.740 2.540 ;
        RECT  6.040 1.700 6.260 2.540 ;
        RECT  3.620 2.080 3.900 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.540 -0.140 7.740 0.600 ;
        RECT  5.890 -0.140 6.170 0.380 ;
        RECT  3.560 -0.140 3.840 0.320 ;
        RECT  1.740 -0.140 1.940 0.640 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.580 0.620 3.020 0.820 ;
        RECT  2.860 1.440 4.180 1.600 ;
        RECT  3.980 1.120 4.180 1.600 ;
        RECT  2.860 0.620 3.020 1.760 ;
        RECT  2.560 1.600 3.020 1.760 ;
        RECT  4.370 0.620 4.580 0.960 ;
        RECT  3.500 0.800 4.580 0.960 ;
        RECT  3.500 0.800 3.700 1.280 ;
        RECT  4.380 0.620 4.580 1.780 ;
        RECT  0.140 0.320 0.340 0.890 ;
        RECT  0.140 0.730 1.020 0.890 ;
        RECT  0.860 0.730 1.020 1.920 ;
        RECT  0.140 1.750 1.020 1.920 ;
        RECT  0.140 1.760 2.270 1.920 ;
        RECT  3.290 1.760 4.220 1.920 ;
        RECT  2.110 1.760 2.270 2.100 ;
        RECT  4.060 1.760 4.220 2.100 ;
        RECT  0.140 1.750 0.340 2.050 ;
        RECT  3.290 1.760 3.450 2.100 ;
        RECT  2.110 1.940 3.450 2.100 ;
        RECT  4.060 1.940 4.730 2.100 ;
        RECT  2.130 0.300 3.340 0.460 ;
        RECT  4.050 0.300 5.500 0.460 ;
        RECT  3.180 0.300 3.340 0.640 ;
        RECT  1.220 0.340 1.580 0.540 ;
        RECT  4.050 0.300 4.210 0.640 ;
        RECT  3.180 0.480 4.210 0.640 ;
        RECT  2.130 0.300 2.300 0.990 ;
        RECT  1.420 0.830 2.300 0.990 ;
        RECT  1.420 0.340 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  5.300 0.300 5.500 1.760 ;
        RECT  5.670 1.160 6.370 1.360 ;
        RECT  4.890 0.620 5.090 2.100 ;
        RECT  5.670 1.160 5.830 2.100 ;
        RECT  4.890 1.940 5.830 2.100 ;
        RECT  5.660 0.680 6.740 0.880 ;
        RECT  6.540 1.100 7.410 1.300 ;
        RECT  6.540 0.370 6.740 1.990 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.730 2.400 ;
        RECT  0.000 1.140 3.730 2.400 ;
        RECT  5.320 1.140 8.000 2.400 ;
        RECT  0.000 1.200 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.730 0.000 8.000 1.140 ;
        RECT  3.730 0.000 5.320 1.200 ;
    END
END DFQM1HM

MACRO DFMQM8HM
    CLASS CORE ;
    FOREIGN DFMQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 4.190 1.300 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.002  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.760 1.440 14.360 1.600 ;
        RECT  14.040 0.310 14.360 1.600 ;
        RECT  13.970 1.440 14.210 2.090 ;
        RECT  12.930 0.690 14.360 0.880 ;
        RECT  13.990 0.310 14.360 0.880 ;
        RECT  12.930 0.350 13.130 0.880 ;
        RECT  12.820 1.440 13.060 2.090 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.510 1.760 14.790 2.540 ;
        RECT  13.360 1.760 13.640 2.540 ;
        RECT  12.240 1.760 12.520 2.540 ;
        RECT  11.120 2.080 11.400 2.540 ;
        RECT  10.120 1.900 10.400 2.540 ;
        RECT  7.080 2.020 7.300 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.590 -0.140 14.790 0.700 ;
        RECT  13.410 -0.140 13.690 0.530 ;
        RECT  12.410 -0.140 12.610 0.620 ;
        RECT  11.390 -0.140 11.610 0.590 ;
        RECT  9.960 -0.140 10.180 0.380 ;
        RECT  7.080 -0.140 7.300 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.580 0.820 ;
        RECT  4.420 1.010 5.040 1.290 ;
        RECT  4.420 0.620 4.580 1.680 ;
        RECT  4.110 1.480 4.580 1.680 ;
        RECT  5.070 0.620 5.380 0.820 ;
        RECT  5.220 0.620 5.380 1.680 ;
        RECT  5.220 0.960 5.690 1.250 ;
        RECT  5.220 0.960 5.420 1.680 ;
        RECT  5.060 1.520 5.420 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.860 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.660 0.300 5.860 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.580 1.660 5.900 2.100 ;
        RECT  3.810 1.940 5.900 2.100 ;
        RECT  6.060 0.320 6.390 0.600 ;
        RECT  6.060 0.320 6.220 1.640 ;
        RECT  7.360 1.180 7.580 1.500 ;
        RECT  6.060 1.340 7.580 1.500 ;
        RECT  6.060 1.340 6.420 1.640 ;
        RECT  6.890 0.860 8.000 1.020 ;
        RECT  6.890 0.860 7.200 1.180 ;
        RECT  7.800 0.620 8.000 1.780 ;
        RECT  7.460 0.300 8.340 0.460 ;
        RECT  7.460 0.300 7.620 0.700 ;
        RECT  6.570 0.540 7.620 0.700 ;
        RECT  8.180 0.300 8.340 1.130 ;
        RECT  6.570 0.540 6.730 1.170 ;
        RECT  6.400 0.890 6.730 1.170 ;
        RECT  6.710 1.700 7.620 1.860 ;
        RECT  7.460 1.700 7.620 2.100 ;
        RECT  6.710 1.700 6.880 2.100 ;
        RECT  6.340 1.900 6.880 2.100 ;
        RECT  7.460 1.940 9.550 2.100 ;
        RECT  9.260 0.620 9.480 1.020 ;
        RECT  10.660 0.620 10.860 1.020 ;
        RECT  9.260 0.860 10.860 1.020 ;
        RECT  9.260 0.620 9.420 1.780 ;
        RECT  9.000 1.500 9.420 1.780 ;
        RECT  9.000 1.560 10.880 1.740 ;
        RECT  9.000 1.560 9.880 1.780 ;
        RECT  10.680 1.560 10.880 1.880 ;
        RECT  8.510 0.300 9.800 0.460 ;
        RECT  10.340 0.300 11.230 0.460 ;
        RECT  9.640 0.300 9.800 0.700 ;
        RECT  8.510 0.300 8.770 0.620 ;
        RECT  10.340 0.300 10.500 0.700 ;
        RECT  9.640 0.540 10.500 0.700 ;
        RECT  11.070 0.300 11.230 1.000 ;
        RECT  11.070 0.840 11.770 1.000 ;
        RECT  11.570 0.840 11.770 1.250 ;
        RECT  8.570 0.300 8.770 1.720 ;
        RECT  8.340 1.490 8.770 1.720 ;
        RECT  11.850 0.410 12.170 0.610 ;
        RECT  11.990 1.050 13.670 1.250 ;
        RECT  9.940 1.180 11.370 1.400 ;
        RECT  11.180 1.180 11.370 1.600 ;
        RECT  11.990 0.410 12.170 1.600 ;
        RECT  11.180 1.440 12.170 1.600 ;
        RECT  11.700 1.440 11.940 2.090 ;
        LAYER VTPH ;
        RECT  11.120 1.080 14.800 2.400 ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.630 1.050 6.830 2.400 ;
        RECT  3.050 1.140 6.830 2.400 ;
        RECT  11.060 1.140 15.200 2.400 ;
        RECT  0.000 1.200 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 1.050 ;
        RECT  6.830 0.000 15.200 1.080 ;
        RECT  0.000 0.000 5.630 1.140 ;
        RECT  6.830 0.000 11.120 1.140 ;
        RECT  14.800 0.000 15.200 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.830 0.000 11.060 1.200 ;
    END
END DFMQM8HM

MACRO DFMQM4HM
    CLASS CORE ;
    FOREIGN DFMQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.452  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.020 0.310 12.190 1.660 ;
        RECT  11.780 1.500 12.080 2.000 ;
        RECT  11.700 0.310 12.190 0.780 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  12.370 1.540 12.590 2.540 ;
        RECT  11.270 1.790 11.550 2.540 ;
        RECT  10.190 1.900 10.470 2.540 ;
        RECT  7.150 2.020 7.370 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  12.350 -0.140 12.550 0.700 ;
        RECT  11.330 -0.140 11.530 0.620 ;
        RECT  10.100 -0.140 10.310 0.680 ;
        RECT  7.150 -0.140 7.370 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.270 0.820 ;
        RECT  4.110 0.620 4.270 1.680 ;
        RECT  4.110 1.010 4.960 1.290 ;
        RECT  4.110 1.010 4.390 1.680 ;
        RECT  4.990 0.620 5.300 0.820 ;
        RECT  5.140 0.620 5.300 1.680 ;
        RECT  5.140 0.960 5.610 1.250 ;
        RECT  5.140 0.960 5.340 1.680 ;
        RECT  4.980 1.480 5.340 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.930 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.730 0.300 5.930 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.650 1.580 5.970 2.100 ;
        RECT  3.810 1.940 5.970 2.100 ;
        RECT  6.130 0.320 6.460 0.600 ;
        RECT  6.130 0.320 6.290 1.640 ;
        RECT  7.430 1.180 7.650 1.500 ;
        RECT  6.130 1.340 7.650 1.500 ;
        RECT  6.130 1.340 6.490 1.640 ;
        RECT  6.960 0.860 8.070 1.020 ;
        RECT  6.960 0.860 7.270 1.180 ;
        RECT  7.870 0.620 8.070 1.780 ;
        RECT  7.530 0.300 8.410 0.460 ;
        RECT  7.530 0.300 7.690 0.700 ;
        RECT  6.640 0.540 7.690 0.700 ;
        RECT  8.250 0.300 8.410 1.130 ;
        RECT  6.640 0.540 6.800 1.170 ;
        RECT  6.470 0.890 6.800 1.170 ;
        RECT  6.780 1.700 7.690 1.860 ;
        RECT  7.530 1.700 7.690 2.100 ;
        RECT  6.780 1.700 6.950 2.100 ;
        RECT  6.410 1.900 6.950 2.100 ;
        RECT  7.530 1.940 9.620 2.100 ;
        RECT  9.330 0.620 9.550 1.780 ;
        RECT  9.070 1.500 9.550 1.780 ;
        RECT  9.070 1.560 9.990 1.780 ;
        RECT  8.580 0.300 9.870 0.460 ;
        RECT  8.580 0.300 8.840 0.620 ;
        RECT  9.710 0.300 9.870 1.000 ;
        RECT  9.710 0.840 10.770 1.000 ;
        RECT  10.570 0.840 10.770 1.250 ;
        RECT  8.640 0.300 8.840 1.720 ;
        RECT  8.410 1.490 8.840 1.720 ;
        RECT  10.750 0.410 11.150 0.610 ;
        RECT  10.930 1.040 11.790 1.250 ;
        RECT  9.770 1.180 10.310 1.400 ;
        RECT  10.150 1.180 10.310 1.660 ;
        RECT  10.930 0.410 11.150 1.660 ;
        RECT  10.150 1.500 11.150 1.660 ;
        RECT  10.740 1.500 11.040 2.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.520 1.050 6.900 2.400 ;
        RECT  3.050 1.140 6.900 2.400 ;
        RECT  9.860 1.140 12.800 2.400 ;
        RECT  0.000 1.200 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.050 ;
        RECT  0.000 0.000 5.520 1.140 ;
        RECT  6.900 0.000 12.800 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.900 0.000 9.860 1.200 ;
    END
END DFMQM4HM

MACRO DFMQM2HM
    CLASS CORE ;
    FOREIGN DFMQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.230 1.460 11.570 2.090 ;
        RECT  11.400 0.440 11.570 2.090 ;
        RECT  11.230 0.440 11.570 0.770 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  11.750 1.400 12.030 2.540 ;
        RECT  10.190 1.900 10.470 2.540 ;
        RECT  7.110 2.020 7.330 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  11.810 -0.140 12.010 0.700 ;
        RECT  10.130 -0.140 10.430 0.630 ;
        RECT  7.110 -0.140 7.330 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.380 0.820 ;
        RECT  4.110 0.620 4.380 1.680 ;
        RECT  4.110 1.010 4.960 1.290 ;
        RECT  4.110 1.010 4.390 1.680 ;
        RECT  4.990 0.620 5.300 0.820 ;
        RECT  5.140 0.620 5.300 1.680 ;
        RECT  5.140 0.960 5.610 1.250 ;
        RECT  5.140 0.960 5.340 1.680 ;
        RECT  4.980 1.480 5.340 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.890 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.690 0.300 5.890 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.610 1.580 5.930 2.100 ;
        RECT  3.810 1.940 5.930 2.100 ;
        RECT  6.090 0.320 6.420 0.600 ;
        RECT  6.090 0.320 6.250 1.640 ;
        RECT  7.390 1.180 7.610 1.500 ;
        RECT  6.090 1.340 7.610 1.500 ;
        RECT  6.090 1.340 6.450 1.640 ;
        RECT  6.920 0.860 8.030 1.020 ;
        RECT  6.920 0.860 7.230 1.180 ;
        RECT  7.830 0.620 8.030 1.780 ;
        RECT  7.490 0.300 8.370 0.460 ;
        RECT  7.490 0.300 7.650 0.700 ;
        RECT  6.600 0.540 7.650 0.700 ;
        RECT  8.210 0.300 8.370 1.130 ;
        RECT  6.600 0.540 6.760 1.170 ;
        RECT  6.430 0.890 6.760 1.170 ;
        RECT  6.740 1.700 7.650 1.860 ;
        RECT  7.490 1.700 7.650 2.100 ;
        RECT  6.740 1.700 6.910 2.100 ;
        RECT  6.370 1.900 6.910 2.100 ;
        RECT  7.490 1.940 9.580 2.100 ;
        RECT  9.290 0.620 9.510 1.780 ;
        RECT  9.030 1.500 9.510 1.780 ;
        RECT  9.030 1.560 9.950 1.780 ;
        RECT  8.540 0.300 9.830 0.460 ;
        RECT  9.670 0.300 9.830 1.000 ;
        RECT  9.670 0.840 10.640 1.000 ;
        RECT  10.430 0.840 10.640 1.250 ;
        RECT  8.540 0.300 8.800 1.720 ;
        RECT  8.370 1.490 8.800 1.720 ;
        RECT  10.810 0.330 11.010 2.090 ;
        RECT  10.810 0.960 11.140 1.240 ;
        RECT  9.730 1.180 10.270 1.380 ;
        RECT  10.110 1.180 10.270 1.660 ;
        RECT  10.110 1.500 11.070 1.660 ;
        RECT  10.810 0.960 11.070 2.090 ;
        RECT  10.720 1.500 11.070 2.090 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.520 1.050 6.860 2.400 ;
        RECT  3.050 1.140 6.860 2.400 ;
        RECT  9.820 1.140 12.400 2.400 ;
        RECT  0.000 1.200 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.050 ;
        RECT  0.000 0.000 5.520 1.140 ;
        RECT  6.860 0.000 12.400 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.860 0.000 9.820 1.200 ;
    END
END DFMQM2HM

MACRO DFMQM1HM
    CLASS CORE ;
    FOREIGN DFMQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.230 1.570 11.550 1.770 ;
        RECT  11.380 0.350 11.550 1.770 ;
        RECT  11.230 0.350 11.550 0.770 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  11.750 1.600 12.030 2.540 ;
        RECT  10.190 1.880 10.470 2.540 ;
        RECT  7.110 2.020 7.330 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  11.810 -0.140 12.010 0.650 ;
        RECT  10.230 -0.140 10.530 0.630 ;
        RECT  7.110 -0.140 7.330 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.380 0.820 ;
        RECT  4.110 0.620 4.380 1.680 ;
        RECT  4.110 1.010 4.960 1.290 ;
        RECT  4.110 1.010 4.390 1.680 ;
        RECT  4.990 0.620 5.300 0.820 ;
        RECT  5.140 0.620 5.300 1.680 ;
        RECT  5.140 0.960 5.610 1.250 ;
        RECT  5.140 0.960 5.340 1.680 ;
        RECT  4.980 1.480 5.340 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.890 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.690 0.300 5.890 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.610 1.560 5.930 2.100 ;
        RECT  3.810 1.940 5.930 2.100 ;
        RECT  6.090 0.320 6.420 0.600 ;
        RECT  6.090 0.320 6.250 1.650 ;
        RECT  7.390 1.180 7.610 1.500 ;
        RECT  6.090 1.340 7.610 1.500 ;
        RECT  6.090 1.340 6.450 1.650 ;
        RECT  6.920 0.860 8.030 1.020 ;
        RECT  6.920 0.860 7.230 1.180 ;
        RECT  7.830 0.620 8.030 1.780 ;
        RECT  7.490 0.300 8.370 0.460 ;
        RECT  7.490 0.300 7.650 0.700 ;
        RECT  6.600 0.540 7.650 0.700 ;
        RECT  8.210 0.300 8.370 1.130 ;
        RECT  6.600 0.540 6.760 1.170 ;
        RECT  6.430 0.890 6.760 1.170 ;
        RECT  6.740 1.700 7.650 1.860 ;
        RECT  7.490 1.700 7.650 2.100 ;
        RECT  6.740 1.700 6.910 2.100 ;
        RECT  6.370 1.900 6.910 2.100 ;
        RECT  7.490 1.940 9.580 2.100 ;
        RECT  9.290 0.620 9.510 1.780 ;
        RECT  9.030 1.500 9.510 1.780 ;
        RECT  9.030 1.560 9.950 1.780 ;
        RECT  8.540 0.300 9.830 0.460 ;
        RECT  9.670 0.300 9.830 1.000 ;
        RECT  9.670 0.840 10.640 1.000 ;
        RECT  10.430 0.840 10.640 1.250 ;
        RECT  8.540 0.300 8.800 1.720 ;
        RECT  8.370 1.490 8.800 1.720 ;
        RECT  10.810 0.330 11.010 1.930 ;
        RECT  10.810 0.960 11.120 1.240 ;
        RECT  9.730 1.180 10.270 1.380 ;
        RECT  10.110 1.180 10.270 1.720 ;
        RECT  10.110 1.560 11.070 1.720 ;
        RECT  10.810 0.960 11.070 1.930 ;
        RECT  10.750 1.560 11.070 1.930 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.520 1.050 6.860 2.400 ;
        RECT  3.050 1.140 6.860 2.400 ;
        RECT  9.820 1.140 12.400 2.400 ;
        RECT  0.000 1.200 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.050 ;
        RECT  0.000 0.000 5.520 1.140 ;
        RECT  6.860 0.000 12.400 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.860 0.000 9.820 1.200 ;
    END
END DFMQM1HM

MACRO DFMM8HM
    CLASS CORE ;
    FOREIGN DFMM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 4.190 1.300 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.002  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.760 1.440 14.360 1.600 ;
        RECT  14.040 0.310 14.360 1.600 ;
        RECT  12.930 0.690 14.360 0.880 ;
        RECT  13.990 0.310 14.360 0.880 ;
        RECT  12.930 0.350 13.130 0.880 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.985  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.150 0.390 16.350 2.100 ;
        RECT  15.110 1.230 16.350 1.560 ;
        RECT  15.110 0.420 15.310 2.100 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 17.200 2.540 ;
        RECT  16.670 1.480 16.870 2.540 ;
        RECT  15.630 1.740 15.830 2.540 ;
        RECT  14.510 2.080 14.790 2.540 ;
        RECT  13.360 2.080 13.640 2.540 ;
        RECT  12.240 2.080 12.520 2.540 ;
        RECT  11.120 2.080 11.400 2.540 ;
        RECT  10.120 1.900 10.400 2.540 ;
        RECT  7.080 2.020 7.300 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 17.200 0.140 ;
        RECT  16.670 -0.140 16.870 0.670 ;
        RECT  15.630 -0.140 15.830 0.670 ;
        RECT  14.590 -0.140 14.790 0.700 ;
        RECT  13.410 -0.140 13.690 0.530 ;
        RECT  12.410 -0.140 12.610 0.620 ;
        RECT  11.390 -0.140 11.610 0.590 ;
        RECT  9.960 -0.140 10.180 0.380 ;
        RECT  7.080 -0.140 7.300 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.580 0.820 ;
        RECT  4.420 1.010 5.040 1.290 ;
        RECT  4.420 0.620 4.580 1.680 ;
        RECT  4.110 1.480 4.580 1.680 ;
        RECT  5.070 0.620 5.380 0.820 ;
        RECT  5.220 0.620 5.380 1.680 ;
        RECT  5.220 0.960 5.690 1.250 ;
        RECT  5.220 0.960 5.420 1.680 ;
        RECT  5.060 1.520 5.420 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.860 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.660 0.300 5.860 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.580 1.660 5.900 2.100 ;
        RECT  3.810 1.940 5.900 2.100 ;
        RECT  6.060 0.320 6.390 0.600 ;
        RECT  6.060 0.320 6.220 1.640 ;
        RECT  7.360 1.180 7.580 1.500 ;
        RECT  6.060 1.340 7.580 1.500 ;
        RECT  6.060 1.340 6.420 1.640 ;
        RECT  6.890 0.860 8.000 1.020 ;
        RECT  6.890 0.860 7.200 1.180 ;
        RECT  7.800 0.620 8.000 1.780 ;
        RECT  7.460 0.300 8.340 0.460 ;
        RECT  7.460 0.300 7.620 0.700 ;
        RECT  6.570 0.540 7.620 0.700 ;
        RECT  8.180 0.300 8.340 1.130 ;
        RECT  6.570 0.540 6.730 1.170 ;
        RECT  6.400 0.890 6.730 1.170 ;
        RECT  6.710 1.700 7.620 1.860 ;
        RECT  7.460 1.700 7.620 2.100 ;
        RECT  6.710 1.700 6.880 2.100 ;
        RECT  6.340 1.900 6.880 2.100 ;
        RECT  7.460 1.940 9.550 2.100 ;
        RECT  8.510 0.300 9.800 0.460 ;
        RECT  10.340 0.300 11.230 0.460 ;
        RECT  9.640 0.300 9.800 0.700 ;
        RECT  8.510 0.300 8.770 0.620 ;
        RECT  10.340 0.300 10.500 0.700 ;
        RECT  9.640 0.540 10.500 0.700 ;
        RECT  11.070 0.300 11.230 1.000 ;
        RECT  11.070 0.840 11.770 1.000 ;
        RECT  11.570 0.840 11.770 1.250 ;
        RECT  8.570 0.300 8.770 1.720 ;
        RECT  8.340 1.490 8.770 1.720 ;
        RECT  11.850 0.410 12.170 0.610 ;
        RECT  11.990 1.050 13.670 1.250 ;
        RECT  9.940 1.180 11.370 1.400 ;
        RECT  11.180 1.180 11.370 1.600 ;
        RECT  11.990 0.410 12.170 1.600 ;
        RECT  11.180 1.440 12.170 1.600 ;
        RECT  9.260 0.620 9.480 1.020 ;
        RECT  10.660 0.620 10.860 1.020 ;
        RECT  9.260 0.860 10.860 1.020 ;
        RECT  9.260 0.620 9.420 1.780 ;
        RECT  9.000 1.500 9.420 1.780 ;
        RECT  9.000 1.560 10.880 1.740 ;
        RECT  10.680 1.560 10.880 1.920 ;
        RECT  9.000 1.560 9.880 1.780 ;
        RECT  14.650 0.930 14.850 1.920 ;
        RECT  10.680 1.760 14.850 1.920 ;
        LAYER VTPH ;
        RECT  11.120 1.080 14.800 2.400 ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.630 1.050 6.830 2.400 ;
        RECT  3.050 1.140 6.830 2.400 ;
        RECT  11.060 1.140 17.200 2.400 ;
        RECT  0.000 1.200 17.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 17.200 1.050 ;
        RECT  6.830 0.000 17.200 1.080 ;
        RECT  0.000 0.000 5.630 1.140 ;
        RECT  6.830 0.000 11.120 1.140 ;
        RECT  14.800 0.000 17.200 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.830 0.000 11.060 1.200 ;
    END
END DFMM8HM

MACRO DFMM4HM
    CLASS CORE ;
    FOREIGN DFMM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.452  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.850 1.440 12.360 1.600 ;
        RECT  12.190 0.310 12.360 1.600 ;
        RECT  11.910 0.310 12.360 0.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.486  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.070 1.200 13.530 1.560 ;
        RECT  13.070 0.420 13.270 2.100 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.590 1.740 13.790 2.540 ;
        RECT  12.470 2.080 12.750 2.540 ;
        RECT  11.350 2.080 11.630 2.540 ;
        RECT  10.230 2.080 10.510 2.540 ;
        RECT  7.150 2.020 7.370 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.590 -0.140 13.790 0.670 ;
        RECT  12.550 -0.140 12.750 0.700 ;
        RECT  11.450 -0.140 11.650 0.620 ;
        RECT  10.170 -0.140 10.470 0.630 ;
        RECT  7.150 -0.140 7.370 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.270 0.820 ;
        RECT  4.110 0.620 4.270 1.680 ;
        RECT  4.110 1.010 4.960 1.290 ;
        RECT  4.110 1.010 4.390 1.680 ;
        RECT  4.990 0.620 5.300 0.820 ;
        RECT  5.140 0.620 5.300 1.680 ;
        RECT  5.140 0.960 5.610 1.250 ;
        RECT  5.140 0.960 5.340 1.680 ;
        RECT  4.980 1.480 5.340 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.930 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.730 0.300 5.930 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.650 1.580 5.970 2.100 ;
        RECT  3.810 1.940 5.970 2.100 ;
        RECT  6.130 0.320 6.460 0.600 ;
        RECT  6.130 0.320 6.290 1.640 ;
        RECT  7.430 1.180 7.650 1.500 ;
        RECT  6.130 1.340 7.650 1.500 ;
        RECT  6.130 1.340 6.490 1.640 ;
        RECT  6.960 0.860 8.070 1.020 ;
        RECT  6.960 0.860 7.270 1.180 ;
        RECT  7.870 0.620 8.070 1.780 ;
        RECT  7.530 0.300 8.410 0.460 ;
        RECT  7.530 0.300 7.690 0.700 ;
        RECT  6.640 0.540 7.690 0.700 ;
        RECT  8.250 0.300 8.410 1.130 ;
        RECT  6.640 0.540 6.800 1.170 ;
        RECT  6.470 0.890 6.800 1.170 ;
        RECT  6.780 1.700 7.690 1.860 ;
        RECT  7.530 1.700 7.690 2.100 ;
        RECT  6.780 1.700 6.950 2.100 ;
        RECT  6.410 1.900 6.950 2.100 ;
        RECT  7.530 1.940 9.620 2.100 ;
        RECT  8.580 0.300 9.870 0.460 ;
        RECT  8.580 0.300 8.840 0.620 ;
        RECT  9.710 0.300 9.870 1.000 ;
        RECT  9.710 0.840 10.950 1.000 ;
        RECT  10.750 0.840 10.950 1.250 ;
        RECT  8.640 0.300 8.840 1.720 ;
        RECT  8.410 1.490 8.840 1.720 ;
        RECT  10.870 0.410 11.290 0.610 ;
        RECT  11.110 1.040 12.010 1.250 ;
        RECT  9.770 1.180 10.310 1.400 ;
        RECT  10.150 1.180 10.310 1.600 ;
        RECT  11.110 0.410 11.290 1.600 ;
        RECT  10.150 1.440 11.290 1.600 ;
        RECT  9.330 0.620 9.550 1.780 ;
        RECT  9.070 1.500 9.550 1.780 ;
        RECT  9.070 1.560 9.990 1.780 ;
        RECT  12.610 0.930 12.810 1.920 ;
        RECT  9.780 1.760 12.810 1.920 ;
        LAYER VTPH ;
        RECT  9.860 1.080 12.760 2.400 ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.520 1.050 6.900 2.400 ;
        RECT  3.050 1.140 6.900 2.400 ;
        RECT  9.860 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.050 ;
        RECT  6.900 0.000 14.000 1.080 ;
        RECT  0.000 0.000 5.520 1.140 ;
        RECT  12.760 0.000 14.000 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.900 0.000 9.860 1.200 ;
    END
END DFMM4HM

MACRO DFMM2HM
    CLASS CORE ;
    FOREIGN DFMM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.142  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.230 1.400 11.730 1.600 ;
        RECT  11.560 0.440 11.730 1.600 ;
        RECT  11.230 0.440 11.730 0.770 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.484  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.390 0.420 12.700 2.100 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.790 2.080 12.070 2.540 ;
        RECT  10.190 2.080 10.470 2.540 ;
        RECT  7.110 2.020 7.330 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.890 -0.140 12.090 0.700 ;
        RECT  10.130 -0.140 10.430 0.630 ;
        RECT  7.110 -0.140 7.330 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.380 0.820 ;
        RECT  4.110 0.620 4.380 1.680 ;
        RECT  4.110 1.010 4.960 1.290 ;
        RECT  4.110 1.010 4.390 1.680 ;
        RECT  4.990 0.620 5.300 0.820 ;
        RECT  5.140 0.620 5.300 1.680 ;
        RECT  5.140 0.960 5.610 1.250 ;
        RECT  5.140 0.960 5.340 1.680 ;
        RECT  4.980 1.480 5.340 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.890 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.690 0.300 5.890 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.610 1.580 5.930 2.100 ;
        RECT  3.810 1.940 5.930 2.100 ;
        RECT  6.090 0.320 6.420 0.600 ;
        RECT  6.090 0.320 6.250 1.640 ;
        RECT  7.390 1.180 7.610 1.500 ;
        RECT  6.090 1.340 7.610 1.500 ;
        RECT  6.090 1.340 6.450 1.640 ;
        RECT  6.920 0.860 8.030 1.020 ;
        RECT  6.920 0.860 7.230 1.180 ;
        RECT  7.830 0.620 8.030 1.780 ;
        RECT  7.490 0.300 8.370 0.460 ;
        RECT  7.490 0.300 7.650 0.700 ;
        RECT  6.600 0.540 7.650 0.700 ;
        RECT  8.210 0.300 8.370 1.130 ;
        RECT  6.600 0.540 6.760 1.170 ;
        RECT  6.430 0.890 6.760 1.170 ;
        RECT  6.740 1.700 7.650 1.860 ;
        RECT  7.490 1.700 7.650 2.100 ;
        RECT  6.740 1.700 6.910 2.100 ;
        RECT  6.370 1.900 6.910 2.100 ;
        RECT  7.490 1.940 9.580 2.100 ;
        RECT  8.540 0.300 9.830 0.460 ;
        RECT  9.670 0.300 9.830 1.000 ;
        RECT  9.670 0.840 10.640 1.000 ;
        RECT  10.430 0.840 10.640 1.250 ;
        RECT  8.540 0.300 8.800 1.720 ;
        RECT  8.370 1.490 8.800 1.720 ;
        RECT  10.810 0.330 11.010 1.600 ;
        RECT  10.810 0.960 11.400 1.240 ;
        RECT  9.730 1.180 10.270 1.380 ;
        RECT  10.110 1.180 10.270 1.600 ;
        RECT  10.810 0.960 11.070 1.600 ;
        RECT  10.110 1.440 11.070 1.600 ;
        RECT  9.290 0.620 9.510 1.780 ;
        RECT  9.030 1.500 9.510 1.780 ;
        RECT  9.030 1.560 9.950 1.780 ;
        RECT  11.930 0.930 12.130 1.920 ;
        RECT  9.740 1.760 12.130 1.920 ;
        LAYER VTPH ;
        RECT  9.820 1.080 12.080 2.400 ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.520 1.050 6.860 2.400 ;
        RECT  3.050 1.140 6.860 2.400 ;
        RECT  9.820 1.140 12.800 2.400 ;
        RECT  0.000 1.200 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.050 ;
        RECT  6.860 0.000 12.800 1.080 ;
        RECT  0.000 0.000 5.520 1.140 ;
        RECT  12.080 0.000 12.800 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.860 0.000 9.820 1.200 ;
    END
END DFMM2HM

MACRO DFMM1HM
    CLASS CORE ;
    FOREIGN DFMM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.980 3.900 1.560 ;
        END
    END CK
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.890 0.820 1.190 1.410 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.050 1.000 3.500 1.560 ;
        END
    END D2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.230 1.400 11.730 1.600 ;
        RECT  11.560 0.350 11.730 1.600 ;
        RECT  11.230 0.350 11.730 0.770 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.357  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.390 0.340 12.700 1.810 ;
        END
    END QB
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 0.790 2.420 1.400 ;
        RECT  1.350 0.790 2.420 0.990 ;
        RECT  1.350 0.480 1.510 0.990 ;
        RECT  0.550 0.480 1.510 0.640 ;
        RECT  0.440 0.700 0.710 1.160 ;
        RECT  0.550 0.480 0.710 1.160 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  11.790 2.080 12.070 2.540 ;
        RECT  10.190 2.080 10.470 2.540 ;
        RECT  7.110 2.020 7.330 2.540 ;
        RECT  3.370 2.080 3.650 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  11.890 -0.140 12.090 0.650 ;
        RECT  10.230 -0.140 10.530 0.630 ;
        RECT  7.110 -0.140 7.330 0.380 ;
        RECT  3.300 -0.140 3.460 0.470 ;
        RECT  0.700 -0.140 0.980 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.310 0.380 0.510 ;
        RECT  0.100 0.310 0.260 2.100 ;
        RECT  1.350 1.230 2.000 1.570 ;
        RECT  0.100 1.570 1.510 1.740 ;
        RECT  0.100 1.570 0.380 2.100 ;
        RECT  2.600 0.620 2.800 1.780 ;
        RECT  2.520 1.580 2.800 1.780 ;
        RECT  3.940 0.620 4.380 0.820 ;
        RECT  4.110 0.620 4.380 1.680 ;
        RECT  4.110 1.010 4.960 1.290 ;
        RECT  4.110 1.010 4.390 1.680 ;
        RECT  4.990 0.620 5.300 0.820 ;
        RECT  5.140 0.620 5.300 1.680 ;
        RECT  5.140 0.960 5.610 1.250 ;
        RECT  5.140 0.960 5.340 1.680 ;
        RECT  4.980 1.480 5.340 1.680 ;
        RECT  1.680 0.300 3.140 0.460 ;
        RECT  3.620 0.300 5.890 0.460 ;
        RECT  1.680 0.300 2.000 0.540 ;
        RECT  5.690 0.300 5.890 0.600 ;
        RECT  2.980 0.300 3.140 0.820 ;
        RECT  3.620 0.300 3.780 0.820 ;
        RECT  2.980 0.660 3.780 0.820 ;
        RECT  3.050 1.760 3.970 1.920 ;
        RECT  1.810 1.820 2.130 2.100 ;
        RECT  3.810 1.760 3.970 2.100 ;
        RECT  3.050 1.760 3.210 2.100 ;
        RECT  1.810 1.940 3.210 2.100 ;
        RECT  5.610 1.560 5.930 2.100 ;
        RECT  3.810 1.940 5.930 2.100 ;
        RECT  6.090 0.320 6.420 0.600 ;
        RECT  6.090 0.320 6.250 1.650 ;
        RECT  7.390 1.180 7.610 1.500 ;
        RECT  6.090 1.340 7.610 1.500 ;
        RECT  6.090 1.340 6.450 1.650 ;
        RECT  6.920 0.860 8.030 1.020 ;
        RECT  6.920 0.860 7.230 1.180 ;
        RECT  7.830 0.620 8.030 1.780 ;
        RECT  7.490 0.300 8.370 0.460 ;
        RECT  7.490 0.300 7.650 0.700 ;
        RECT  6.600 0.540 7.650 0.700 ;
        RECT  8.210 0.300 8.370 1.130 ;
        RECT  6.600 0.540 6.760 1.170 ;
        RECT  6.430 0.890 6.760 1.170 ;
        RECT  6.740 1.700 7.650 1.860 ;
        RECT  7.490 1.700 7.650 2.100 ;
        RECT  6.740 1.700 6.910 2.100 ;
        RECT  6.370 1.900 6.910 2.100 ;
        RECT  7.490 1.940 9.580 2.100 ;
        RECT  8.540 0.300 9.830 0.460 ;
        RECT  9.670 0.300 9.830 1.000 ;
        RECT  9.670 0.840 10.640 1.000 ;
        RECT  10.430 0.840 10.640 1.250 ;
        RECT  8.540 0.300 8.800 1.720 ;
        RECT  8.370 1.490 8.800 1.720 ;
        RECT  10.810 0.330 11.010 1.600 ;
        RECT  10.810 0.960 11.400 1.240 ;
        RECT  9.730 1.180 10.270 1.380 ;
        RECT  10.110 1.180 10.270 1.600 ;
        RECT  10.810 0.960 11.070 1.600 ;
        RECT  10.110 1.440 11.070 1.600 ;
        RECT  9.290 0.620 9.510 1.780 ;
        RECT  9.030 1.500 9.510 1.780 ;
        RECT  9.030 1.560 9.950 1.780 ;
        RECT  11.930 0.930 12.130 1.920 ;
        RECT  9.740 1.760 12.130 1.920 ;
        LAYER VTPH ;
        RECT  9.820 1.080 12.080 2.400 ;
        RECT  0.000 1.140 2.370 2.400 ;
        RECT  5.520 1.050 6.860 2.400 ;
        RECT  3.050 1.140 6.860 2.400 ;
        RECT  9.820 1.140 12.800 2.400 ;
        RECT  0.000 1.200 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.050 ;
        RECT  6.860 0.000 12.800 1.080 ;
        RECT  0.000 0.000 5.520 1.140 ;
        RECT  12.080 0.000 12.800 1.140 ;
        RECT  2.370 0.000 3.050 1.200 ;
        RECT  6.860 0.000 9.820 1.200 ;
    END
END DFMM1HM

MACRO DFM8HM
    CLASS CORE ;
    FOREIGN DFM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.050 0.590 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.240 2.710 1.460 ;
        RECT  2.430 1.120 2.710 1.460 ;
        RECT  2.040 1.240 2.370 1.500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.412  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.750 1.130 11.040 2.100 ;
        RECT  10.760 0.620 11.040 2.100 ;
        RECT  9.360 1.130 11.040 1.320 ;
        RECT  9.690 1.130 9.940 2.100 ;
        RECT  9.360 0.620 9.640 1.320 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.000 1.220 13.310 2.060 ;
        RECT  13.010 0.430 13.310 2.060 ;
        RECT  11.970 1.220 13.310 1.560 ;
        RECT  11.970 0.440 12.260 2.060 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.540 1.530 13.820 2.540 ;
        RECT  12.560 1.800 12.720 2.540 ;
        RECT  11.450 1.520 11.740 2.540 ;
        RECT  10.210 1.820 10.410 2.540 ;
        RECT  9.050 1.480 9.250 2.540 ;
        RECT  8.010 1.800 8.210 2.540 ;
        RECT  6.860 1.900 7.150 2.540 ;
        RECT  3.690 2.080 3.970 2.540 ;
        RECT  1.630 2.080 1.910 2.540 ;
        RECT  0.670 2.080 0.950 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.540 -0.140 13.800 0.750 ;
        RECT  12.520 -0.140 12.760 0.730 ;
        RECT  11.520 -0.140 11.760 0.740 ;
        RECT  10.120 -0.140 10.280 0.650 ;
        RECT  8.620 -0.140 8.870 0.630 ;
        RECT  7.630 -0.140 7.840 0.600 ;
        RECT  6.170 -0.140 6.380 0.630 ;
        RECT  3.690 -0.140 3.970 0.320 ;
        RECT  1.750 -0.140 1.950 0.640 ;
        RECT  0.630 -0.140 0.910 0.550 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.650 0.620 3.030 0.820 ;
        RECT  3.950 1.170 4.230 1.600 ;
        RECT  2.870 1.440 4.230 1.600 ;
        RECT  2.870 0.620 3.030 1.780 ;
        RECT  2.570 1.620 3.030 1.780 ;
        RECT  3.470 0.800 4.650 0.960 ;
        RECT  3.470 0.800 3.750 1.280 ;
        RECT  4.450 0.620 4.650 1.780 ;
        RECT  0.150 0.440 0.350 0.890 ;
        RECT  0.150 0.730 1.030 0.890 ;
        RECT  0.870 0.730 1.030 1.920 ;
        RECT  0.110 1.720 1.030 1.920 ;
        RECT  0.110 1.760 2.280 1.920 ;
        RECT  3.300 1.760 4.290 1.920 ;
        RECT  2.120 1.760 2.280 2.100 ;
        RECT  4.130 1.760 4.290 2.100 ;
        RECT  3.300 1.760 3.460 2.100 ;
        RECT  2.120 1.940 3.460 2.100 ;
        RECT  4.130 1.940 4.920 2.100 ;
        RECT  2.140 0.300 3.460 0.460 ;
        RECT  4.130 0.300 5.150 0.460 ;
        RECT  3.300 0.300 3.460 0.640 ;
        RECT  4.130 0.300 4.290 0.640 ;
        RECT  3.300 0.480 4.290 0.640 ;
        RECT  1.230 0.450 1.590 0.650 ;
        RECT  2.140 0.300 2.310 0.990 ;
        RECT  1.430 0.830 2.310 0.990 ;
        RECT  1.430 0.450 1.590 1.600 ;
        RECT  1.240 1.400 1.590 1.600 ;
        RECT  4.910 0.680 5.240 0.880 ;
        RECT  6.040 1.110 6.710 1.270 ;
        RECT  5.080 0.680 5.240 2.100 ;
        RECT  6.040 1.110 6.200 2.100 ;
        RECT  5.080 1.940 6.200 2.100 ;
        RECT  6.870 0.620 7.150 1.280 ;
        RECT  6.870 1.120 8.530 1.280 ;
        RECT  6.870 0.620 7.110 1.740 ;
        RECT  6.360 1.580 7.660 1.740 ;
        RECT  6.360 1.580 6.560 2.100 ;
        RECT  7.460 1.580 7.660 2.100 ;
        RECT  6.540 0.300 7.470 0.460 ;
        RECT  9.040 0.300 9.960 0.460 ;
        RECT  10.440 0.300 11.360 0.460 ;
        RECT  5.620 0.620 5.840 1.780 ;
        RECT  8.110 0.320 8.340 0.960 ;
        RECT  7.310 0.300 7.470 0.960 ;
        RECT  8.110 0.790 9.200 0.960 ;
        RECT  9.800 0.300 9.960 0.970 ;
        RECT  6.540 0.300 6.710 0.950 ;
        RECT  5.620 0.790 6.710 0.950 ;
        RECT  9.040 0.300 9.200 0.960 ;
        RECT  7.310 0.800 9.200 0.960 ;
        RECT  10.440 0.300 10.600 0.970 ;
        RECT  9.800 0.810 10.600 0.970 ;
        RECT  11.200 0.300 11.360 1.320 ;
        RECT  11.200 1.030 11.790 1.320 ;
        RECT  5.620 0.790 5.860 1.780 ;
        RECT  8.690 0.790 8.850 2.100 ;
        RECT  8.490 1.500 8.850 2.100 ;
        LAYER VTPH ;
        RECT  1.000 1.080 1.740 2.400 ;
        RECT  0.000 1.140 3.740 2.400 ;
        RECT  6.060 1.140 14.000 2.400 ;
        RECT  0.000 1.200 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 1.000 1.140 ;
        RECT  1.740 0.000 14.000 1.140 ;
        RECT  3.740 0.000 6.060 1.200 ;
    END
END DFM8HM

MACRO DFM4HM
    CLASS CORE ;
    FOREIGN DFM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.050 0.580 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.240 2.700 1.460 ;
        RECT  2.420 1.120 2.700 1.460 ;
        RECT  2.040 1.240 2.360 1.500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.813  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.440 1.620 8.960 2.100 ;
        RECT  8.680 0.620 8.960 2.100 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.890 1.200 10.700 1.560 ;
        RECT  9.890 0.440 10.180 2.060 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.800 2.540 ;
        RECT  10.480 1.800 10.640 2.540 ;
        RECT  9.370 1.520 9.660 2.540 ;
        RECT  8.010 1.810 8.210 2.540 ;
        RECT  6.930 1.840 7.130 2.540 ;
        RECT  3.680 2.080 3.960 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.800 0.140 ;
        RECT  10.460 -0.140 10.680 0.730 ;
        RECT  9.440 -0.140 9.680 0.740 ;
        RECT  8.040 -0.140 8.200 0.630 ;
        RECT  7.100 -0.140 7.300 0.400 ;
        RECT  3.680 -0.140 3.960 0.320 ;
        RECT  1.740 -0.140 1.940 0.640 ;
        RECT  0.620 -0.140 0.900 0.550 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.640 0.620 3.020 0.820 ;
        RECT  3.940 1.170 4.220 1.600 ;
        RECT  2.860 1.440 4.220 1.600 ;
        RECT  2.860 0.620 3.020 1.780 ;
        RECT  2.560 1.620 3.020 1.780 ;
        RECT  3.460 0.800 4.640 0.960 ;
        RECT  3.460 0.800 3.740 1.280 ;
        RECT  4.440 0.620 4.640 1.780 ;
        RECT  0.140 0.330 0.340 0.890 ;
        RECT  0.140 0.730 1.020 0.890 ;
        RECT  0.860 0.730 1.020 1.920 ;
        RECT  0.100 1.750 1.020 1.920 ;
        RECT  0.100 1.760 2.270 1.920 ;
        RECT  3.290 1.760 4.280 1.920 ;
        RECT  2.110 1.760 2.270 2.100 ;
        RECT  4.120 1.760 4.280 2.100 ;
        RECT  0.100 1.750 0.400 2.010 ;
        RECT  3.290 1.760 3.450 2.100 ;
        RECT  2.110 1.940 3.450 2.100 ;
        RECT  4.120 1.940 4.910 2.100 ;
        RECT  2.130 0.300 3.450 0.460 ;
        RECT  4.120 0.300 5.140 0.460 ;
        RECT  3.290 0.300 3.450 0.640 ;
        RECT  1.220 0.340 1.580 0.540 ;
        RECT  4.120 0.300 4.280 0.640 ;
        RECT  3.290 0.480 4.280 0.640 ;
        RECT  2.130 0.300 2.300 0.990 ;
        RECT  1.420 0.830 2.300 0.990 ;
        RECT  1.420 0.340 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  4.900 0.680 5.230 0.880 ;
        RECT  6.030 1.200 6.740 1.360 ;
        RECT  5.070 0.680 5.230 2.100 ;
        RECT  6.030 1.200 6.210 2.100 ;
        RECT  5.070 1.940 6.210 2.100 ;
        RECT  6.300 0.620 6.580 1.040 ;
        RECT  6.300 0.880 7.190 1.040 ;
        RECT  7.030 1.120 7.900 1.280 ;
        RECT  7.030 0.880 7.190 1.680 ;
        RECT  6.430 1.520 7.190 1.680 ;
        RECT  6.430 1.520 6.630 2.100 ;
        RECT  5.610 0.300 6.940 0.460 ;
        RECT  8.360 0.300 9.280 0.460 ;
        RECT  6.780 0.300 6.940 0.720 ;
        RECT  6.780 0.560 7.710 0.720 ;
        RECT  7.480 0.560 7.710 0.960 ;
        RECT  8.360 0.300 8.520 0.950 ;
        RECT  7.480 0.790 8.520 0.950 ;
        RECT  7.480 0.790 8.220 0.960 ;
        RECT  9.120 0.300 9.280 1.320 ;
        RECT  9.120 1.030 9.710 1.320 ;
        RECT  8.060 0.790 8.220 1.600 ;
        RECT  7.450 1.440 8.220 1.600 ;
        RECT  5.610 0.300 5.850 1.780 ;
        RECT  7.450 1.440 7.670 2.100 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.730 2.400 ;
        RECT  0.000 1.140 3.730 2.400 ;
        RECT  6.050 1.140 10.800 2.400 ;
        RECT  0.000 1.200 10.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.800 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.730 0.000 10.800 1.140 ;
        RECT  3.730 0.000 6.050 1.200 ;
    END
END DFM4HM

MACRO DFM2HM
    CLASS CORE ;
    FOREIGN DFM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.050 0.580 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.240 2.700 1.400 ;
        RECT  2.420 1.120 2.700 1.400 ;
        RECT  2.040 1.240 2.360 1.500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.522  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.440 1.440 8.960 2.100 ;
        RECT  8.680 0.620 8.960 2.100 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.890 1.180 10.300 1.610 ;
        RECT  9.890 1.180 10.180 2.060 ;
        RECT  9.890 0.440 10.120 2.060 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.370 1.520 9.660 2.540 ;
        RECT  8.010 1.810 8.210 2.540 ;
        RECT  6.930 1.840 7.130 2.540 ;
        RECT  3.680 2.080 3.960 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.440 -0.140 9.680 0.740 ;
        RECT  8.040 -0.140 8.200 0.630 ;
        RECT  6.950 -0.140 7.150 0.400 ;
        RECT  3.680 -0.140 3.960 0.320 ;
        RECT  1.740 -0.140 1.940 0.640 ;
        RECT  0.620 -0.140 0.900 0.550 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.640 0.620 3.020 0.820 ;
        RECT  2.860 1.440 4.220 1.600 ;
        RECT  3.940 1.170 4.220 1.600 ;
        RECT  2.860 0.620 3.020 1.760 ;
        RECT  2.560 1.600 3.020 1.760 ;
        RECT  3.460 0.800 4.640 0.960 ;
        RECT  3.460 0.800 3.740 1.280 ;
        RECT  4.440 0.620 4.640 1.780 ;
        RECT  0.140 0.330 0.340 0.890 ;
        RECT  0.140 0.730 1.020 0.890 ;
        RECT  0.860 0.730 1.020 1.920 ;
        RECT  0.100 1.750 1.020 1.920 ;
        RECT  0.100 1.760 2.270 1.920 ;
        RECT  3.290 1.760 4.280 1.920 ;
        RECT  2.110 1.760 2.270 2.100 ;
        RECT  4.120 1.760 4.280 2.100 ;
        RECT  0.100 1.750 0.400 2.010 ;
        RECT  3.290 1.760 3.450 2.100 ;
        RECT  2.110 1.940 3.450 2.100 ;
        RECT  4.120 1.940 4.910 2.100 ;
        RECT  2.130 0.300 3.450 0.460 ;
        RECT  4.120 0.300 5.140 0.460 ;
        RECT  3.290 0.300 3.450 0.640 ;
        RECT  1.220 0.340 1.580 0.540 ;
        RECT  4.120 0.300 4.280 0.640 ;
        RECT  3.290 0.480 4.280 0.640 ;
        RECT  2.130 0.300 2.300 0.990 ;
        RECT  1.420 0.830 2.300 0.990 ;
        RECT  1.420 0.340 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  4.900 0.680 5.230 0.880 ;
        RECT  6.030 1.200 6.740 1.360 ;
        RECT  5.070 0.680 5.230 2.100 ;
        RECT  6.030 1.200 6.210 2.100 ;
        RECT  5.070 1.940 6.210 2.100 ;
        RECT  6.150 0.620 6.430 1.040 ;
        RECT  6.150 0.880 7.190 1.040 ;
        RECT  7.030 1.120 7.900 1.280 ;
        RECT  7.030 0.880 7.190 1.680 ;
        RECT  6.430 1.520 7.190 1.680 ;
        RECT  6.430 1.520 6.630 2.100 ;
        RECT  5.610 0.300 6.790 0.460 ;
        RECT  8.360 0.300 9.280 0.460 ;
        RECT  6.630 0.300 6.790 0.720 ;
        RECT  6.630 0.560 7.710 0.720 ;
        RECT  7.370 0.560 7.710 0.960 ;
        RECT  8.360 0.300 8.520 0.950 ;
        RECT  7.370 0.790 8.520 0.950 ;
        RECT  7.370 0.790 8.220 0.960 ;
        RECT  9.120 0.300 9.280 1.320 ;
        RECT  9.120 1.030 9.710 1.320 ;
        RECT  8.060 0.790 8.220 1.600 ;
        RECT  7.390 1.440 8.220 1.600 ;
        RECT  7.390 1.440 7.610 1.760 ;
        RECT  5.610 0.300 5.850 1.780 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.730 2.400 ;
        RECT  0.000 1.140 3.730 2.400 ;
        RECT  6.050 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.730 0.000 10.400 1.140 ;
        RECT  3.730 0.000 6.050 1.200 ;
    END
END DFM2HM

MACRO DFM1HM
    CLASS CORE ;
    FOREIGN DFM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.050 0.580 1.560 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 1.240 2.700 1.400 ;
        RECT  2.420 1.120 2.700 1.400 ;
        RECT  2.040 1.240 2.360 1.500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.414  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.680 0.620 8.960 0.840 ;
        RECT  8.440 1.640 8.840 2.100 ;
        RECT  8.680 0.620 8.840 2.100 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.890 1.170 10.300 1.610 ;
        RECT  9.890 0.420 10.180 2.060 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.380 1.790 9.660 2.540 ;
        RECT  8.010 1.810 8.210 2.540 ;
        RECT  6.930 1.840 7.130 2.540 ;
        RECT  3.680 2.080 3.960 2.540 ;
        RECT  1.620 2.080 1.900 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.440 -0.140 9.680 0.670 ;
        RECT  8.040 -0.140 8.200 0.630 ;
        RECT  6.950 -0.140 7.150 0.400 ;
        RECT  3.680 -0.140 3.960 0.320 ;
        RECT  1.740 -0.140 1.940 0.640 ;
        RECT  0.620 -0.140 0.900 0.550 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.640 0.620 3.020 0.820 ;
        RECT  2.860 1.440 4.220 1.600 ;
        RECT  3.940 1.170 4.220 1.600 ;
        RECT  2.860 0.620 3.020 1.760 ;
        RECT  2.560 1.600 3.020 1.760 ;
        RECT  3.460 0.800 4.640 0.960 ;
        RECT  3.460 0.800 3.740 1.280 ;
        RECT  4.440 0.620 4.640 1.780 ;
        RECT  0.140 0.330 0.340 0.890 ;
        RECT  0.140 0.730 1.020 0.890 ;
        RECT  0.860 0.730 1.020 1.920 ;
        RECT  0.100 1.750 1.020 1.920 ;
        RECT  0.100 1.760 2.270 1.920 ;
        RECT  3.290 1.760 4.280 1.920 ;
        RECT  2.110 1.760 2.270 2.100 ;
        RECT  4.120 1.760 4.280 2.100 ;
        RECT  0.100 1.750 0.400 1.990 ;
        RECT  3.290 1.760 3.450 2.100 ;
        RECT  2.110 1.940 3.450 2.100 ;
        RECT  4.120 1.940 4.910 2.100 ;
        RECT  2.130 0.300 3.450 0.460 ;
        RECT  4.120 0.300 5.140 0.460 ;
        RECT  3.290 0.300 3.450 0.640 ;
        RECT  1.220 0.340 1.580 0.550 ;
        RECT  4.120 0.300 4.280 0.640 ;
        RECT  3.290 0.480 4.280 0.640 ;
        RECT  2.130 0.300 2.300 0.990 ;
        RECT  1.420 0.830 2.300 0.990 ;
        RECT  1.420 0.340 1.580 1.600 ;
        RECT  1.230 1.400 1.580 1.600 ;
        RECT  4.900 0.680 5.230 0.880 ;
        RECT  6.030 1.200 6.740 1.360 ;
        RECT  5.070 0.680 5.230 2.100 ;
        RECT  6.030 1.200 6.210 2.100 ;
        RECT  5.070 1.940 6.210 2.100 ;
        RECT  6.150 0.620 6.430 1.040 ;
        RECT  6.150 0.880 7.190 1.040 ;
        RECT  7.030 1.120 7.900 1.280 ;
        RECT  7.030 0.880 7.190 1.680 ;
        RECT  6.430 1.520 7.190 1.680 ;
        RECT  6.430 1.520 6.630 2.100 ;
        RECT  5.610 0.300 6.790 0.460 ;
        RECT  8.360 0.300 9.280 0.460 ;
        RECT  6.630 0.300 6.790 0.720 ;
        RECT  6.630 0.560 7.710 0.720 ;
        RECT  7.370 0.560 7.710 0.960 ;
        RECT  8.360 0.300 8.520 0.950 ;
        RECT  7.370 0.790 8.520 0.950 ;
        RECT  7.370 0.790 8.220 0.960 ;
        RECT  9.120 0.300 9.280 1.320 ;
        RECT  9.120 1.030 9.710 1.320 ;
        RECT  8.060 0.790 8.220 1.600 ;
        RECT  7.390 1.440 8.220 1.600 ;
        RECT  7.390 1.440 7.610 1.760 ;
        RECT  5.610 0.300 5.850 1.780 ;
        LAYER VTPH ;
        RECT  0.990 1.080 1.730 2.400 ;
        RECT  0.000 1.140 3.730 2.400 ;
        RECT  6.050 1.140 10.400 2.400 ;
        RECT  0.000 1.200 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 0.990 1.140 ;
        RECT  1.730 0.000 10.400 1.140 ;
        RECT  3.730 0.000 6.050 1.200 ;
    END
END DFM1HM

MACRO DFEZRM8HM
    CLASS CORE ;
    FOREIGN DFEZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.104  LAYER ME1  ;
        ANTENNAGATEAREA 0.104  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.586  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.060 3.500 1.260 ;
        LAYER ME2 ;
        RECT  3.300 0.810 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.120 1.040 3.600 1.280 ;
        END
    END RB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.036  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.950 1.900 1.150 ;
        LAYER ME2 ;
        RECT  1.700 0.700 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.500 0.950 2.080 1.230 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        ANTENNAGATEAREA 0.220  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.871  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 0.950 0.700 1.150 ;
        LAYER ME2 ;
        RECT  0.500 0.700 0.700 1.340 ;
        LAYER ME1 ;
        RECT  0.500 0.810 0.760 1.340 ;
        END
    END E
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.240 0.840 4.860 1.190 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.888  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.860 1.400 17.350 1.600 ;
        RECT  17.040 0.400 17.350 1.600 ;
        RECT  16.080 1.250 17.350 1.600 ;
        RECT  16.080 0.400 16.280 1.600 ;
        RECT  15.990 0.400 16.280 0.680 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.980  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  19.140 0.400 19.500 2.100 ;
        RECT  18.080 0.840 19.500 1.150 ;
        RECT  18.080 0.840 18.400 2.060 ;
        RECT  18.080 0.400 18.390 2.060 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 20.000 2.540 ;
        RECT  19.660 1.480 19.860 2.540 ;
        RECT  18.620 1.470 18.820 2.540 ;
        RECT  16.460 2.080 16.740 2.540 ;
        RECT  15.300 2.080 15.580 2.540 ;
        RECT  14.180 2.080 14.460 2.540 ;
        RECT  12.960 1.900 13.240 2.540 ;
        RECT  8.440 1.860 8.720 2.540 ;
        RECT  4.450 1.860 4.730 2.540 ;
        RECT  2.680 2.080 2.960 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 20.000 0.140 ;
        RECT  19.660 -0.140 19.860 0.680 ;
        RECT  18.620 -0.140 18.820 0.680 ;
        RECT  17.580 -0.140 17.780 0.680 ;
        RECT  16.520 -0.140 16.760 0.680 ;
        RECT  15.500 -0.140 15.700 0.680 ;
        RECT  14.480 -0.140 14.640 0.680 ;
        RECT  12.960 -0.140 13.240 0.320 ;
        RECT  8.900 -0.140 9.180 0.540 ;
        RECT  3.480 -0.140 3.700 0.410 ;
        RECT  0.620 -0.140 0.900 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.960 1.440 2.460 1.600 ;
        RECT  2.260 0.940 2.460 1.600 ;
        RECT  0.960 0.910 1.160 1.660 ;
        RECT  0.140 1.500 1.160 1.660 ;
        RECT  0.140 0.410 0.340 2.030 ;
        RECT  1.100 0.300 3.240 0.460 ;
        RECT  2.920 0.300 3.240 0.560 ;
        RECT  1.100 0.300 1.380 0.590 ;
        RECT  2.760 1.160 2.960 1.600 ;
        RECT  3.770 1.040 3.970 1.600 ;
        RECT  2.760 1.440 3.970 1.600 ;
        RECT  5.160 0.620 5.440 0.840 ;
        RECT  5.210 0.620 5.440 1.760 ;
        RECT  5.210 0.970 6.080 1.250 ;
        RECT  5.210 0.970 5.480 1.760 ;
        RECT  6.200 0.620 6.540 0.820 ;
        RECT  6.240 0.620 6.540 1.220 ;
        RECT  6.240 0.930 6.580 1.220 ;
        RECT  6.240 0.620 6.520 1.730 ;
        RECT  3.860 0.300 6.920 0.460 ;
        RECT  6.720 0.300 6.920 0.600 ;
        RECT  1.880 0.620 2.770 0.780 ;
        RECT  3.860 0.300 4.020 0.880 ;
        RECT  2.610 0.720 4.020 0.880 ;
        RECT  4.130 1.540 5.050 1.700 ;
        RECT  4.130 1.540 4.290 1.920 ;
        RECT  1.660 1.760 4.290 1.920 ;
        RECT  4.890 1.540 5.050 2.100 ;
        RECT  1.660 1.760 1.860 2.080 ;
        RECT  6.720 1.480 6.950 2.100 ;
        RECT  4.890 1.940 6.950 2.100 ;
        RECT  7.390 0.370 7.700 0.710 ;
        RECT  7.390 0.370 7.590 1.650 ;
        RECT  7.390 1.340 9.220 1.500 ;
        RECT  7.390 1.340 7.840 1.650 ;
        RECT  9.000 1.340 9.220 1.840 ;
        RECT  8.600 1.020 9.970 1.180 ;
        RECT  9.690 0.660 9.970 1.800 ;
        RECT  9.680 1.020 9.970 1.800 ;
        RECT  9.680 1.480 10.040 1.800 ;
        RECT  9.360 0.300 10.380 0.460 ;
        RECT  9.360 0.300 9.530 0.860 ;
        RECT  7.980 0.700 9.530 0.860 ;
        RECT  7.980 0.700 8.180 1.180 ;
        RECT  10.180 0.300 10.380 1.180 ;
        RECT  10.670 0.300 12.800 0.460 ;
        RECT  13.400 0.300 14.320 0.460 ;
        RECT  12.620 0.300 12.800 0.660 ;
        RECT  13.400 0.300 13.560 0.660 ;
        RECT  12.620 0.500 13.560 0.660 ;
        RECT  14.160 0.300 14.320 1.270 ;
        RECT  10.670 0.300 10.940 1.780 ;
        RECT  14.980 0.950 15.900 1.230 ;
        RECT  12.600 1.160 13.920 1.360 ;
        RECT  13.760 1.160 13.920 1.600 ;
        RECT  14.980 0.400 15.180 1.600 ;
        RECT  13.760 1.440 15.180 1.600 ;
        RECT  12.180 0.620 12.460 1.000 ;
        RECT  13.720 0.620 14.000 1.000 ;
        RECT  12.180 0.840 14.000 1.000 ;
        RECT  11.370 1.330 12.370 1.610 ;
        RECT  12.070 1.540 13.600 1.700 ;
        RECT  13.430 1.540 13.600 1.920 ;
        RECT  17.720 0.940 17.920 1.920 ;
        RECT  13.430 1.760 17.920 1.920 ;
        RECT  12.180 0.620 12.370 2.100 ;
        RECT  12.070 1.330 12.370 2.100 ;
        LAYER VTPH ;
        RECT  6.760 0.970 7.880 2.400 ;
        RECT  0.420 1.040 1.750 2.400 ;
        RECT  10.690 1.020 11.910 2.400 ;
        RECT  10.240 1.090 11.910 2.400 ;
        RECT  14.180 1.080 19.460 2.400 ;
        RECT  6.760 1.060 8.580 2.400 ;
        RECT  0.000 1.140 8.580 2.400 ;
        RECT  10.240 1.140 20.000 2.400 ;
        RECT  0.000 1.180 20.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 20.000 0.970 ;
        RECT  7.880 0.000 20.000 1.020 ;
        RECT  0.000 0.000 6.760 1.040 ;
        RECT  7.880 0.000 10.690 1.060 ;
        RECT  11.910 0.000 20.000 1.080 ;
        RECT  8.580 0.000 10.690 1.090 ;
        RECT  0.000 0.000 0.420 1.140 ;
        RECT  1.750 0.000 6.760 1.140 ;
        RECT  11.910 0.000 14.180 1.140 ;
        RECT  19.460 0.000 20.000 1.140 ;
        RECT  8.580 0.000 10.240 1.180 ;
    END
END DFEZRM8HM

MACRO DFEZRM4HM
    CLASS CORE ;
    FOREIGN DFEZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.036  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.950 1.900 1.150 ;
        LAYER ME2 ;
        RECT  1.700 0.700 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.500 0.950 2.080 1.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        ANTENNAGATEAREA 0.059  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.898  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.180 1.050 4.380 1.250 ;
        LAYER ME2 ;
        RECT  4.100 0.810 4.380 1.610 ;
        LAYER ME1 ;
        RECT  4.180 0.940 4.540 1.360 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.540  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.170 1.400 14.700 1.600 ;
        RECT  14.390 0.400 14.700 1.600 ;
        RECT  14.180 0.400 14.700 0.680 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.300 1.440 16.300 1.600 ;
        RECT  16.040 0.720 16.300 1.600 ;
        RECT  15.300 0.720 16.300 0.880 ;
        RECT  15.300 1.440 15.590 2.100 ;
        RECT  15.300 0.400 15.590 0.880 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        ANTENNAGATEAREA 0.220  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.729  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 0.950 0.700 1.150 ;
        LAYER ME2 ;
        RECT  0.500 0.700 0.700 1.340 ;
        LAYER ME1 ;
        RECT  0.500 0.810 0.760 1.280 ;
        END
    END E
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.486  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.220 1.260 3.420 1.460 ;
        LAYER ME2 ;
        RECT  3.220 0.810 3.500 1.610 ;
        LAYER ME1 ;
        RECT  3.120 1.260 3.520 1.600 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.400 2.540 ;
        RECT  15.930 1.790 16.130 2.540 ;
        RECT  14.810 2.080 15.090 2.540 ;
        RECT  13.610 2.080 13.890 2.540 ;
        RECT  12.450 2.080 12.730 2.540 ;
        RECT  7.930 1.860 8.210 2.540 ;
        RECT  4.070 1.860 4.350 2.540 ;
        RECT  2.680 2.080 2.960 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.400 0.140 ;
        RECT  15.930 -0.140 16.130 0.560 ;
        RECT  14.910 -0.140 15.110 0.720 ;
        RECT  13.610 -0.140 13.810 0.680 ;
        RECT  12.550 -0.140 12.710 0.600 ;
        RECT  8.390 -0.140 8.670 0.540 ;
        RECT  3.580 -0.140 3.800 0.410 ;
        RECT  0.620 -0.140 0.900 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.960 0.910 1.160 1.600 ;
        RECT  2.260 0.940 2.460 1.600 ;
        RECT  0.140 1.440 2.460 1.600 ;
        RECT  0.140 0.410 0.340 2.030 ;
        RECT  1.100 0.300 3.310 0.460 ;
        RECT  1.100 0.300 1.380 0.590 ;
        RECT  2.760 0.940 3.990 1.100 ;
        RECT  3.770 0.940 3.990 1.340 ;
        RECT  2.760 0.940 2.960 1.500 ;
        RECT  4.770 0.620 5.060 0.840 ;
        RECT  4.830 0.620 5.060 1.760 ;
        RECT  4.830 0.970 5.570 1.250 ;
        RECT  4.830 0.970 5.100 1.760 ;
        RECT  5.690 0.620 6.030 0.820 ;
        RECT  5.730 0.620 6.030 1.220 ;
        RECT  5.730 0.930 6.070 1.220 ;
        RECT  5.730 0.620 6.010 1.730 ;
        RECT  3.960 0.300 6.410 0.460 ;
        RECT  6.210 0.300 6.410 0.600 ;
        RECT  3.960 0.300 4.120 0.780 ;
        RECT  1.880 0.620 4.120 0.780 ;
        RECT  3.750 1.540 4.670 1.700 ;
        RECT  3.750 1.540 3.910 1.920 ;
        RECT  1.660 1.760 3.910 1.920 ;
        RECT  4.510 1.540 4.670 2.100 ;
        RECT  1.660 1.760 1.860 2.080 ;
        RECT  6.210 1.480 6.440 2.100 ;
        RECT  4.510 1.940 6.440 2.100 ;
        RECT  6.880 0.370 7.190 0.710 ;
        RECT  6.880 0.370 7.080 1.650 ;
        RECT  6.880 1.340 8.710 1.500 ;
        RECT  6.880 1.340 7.330 1.650 ;
        RECT  8.490 1.340 8.710 1.840 ;
        RECT  8.090 1.020 9.460 1.180 ;
        RECT  9.180 0.660 9.460 1.800 ;
        RECT  9.170 1.020 9.460 1.800 ;
        RECT  9.170 1.480 9.530 1.800 ;
        RECT  8.850 0.300 9.870 0.460 ;
        RECT  8.850 0.300 9.020 0.860 ;
        RECT  7.470 0.700 9.020 0.860 ;
        RECT  7.470 0.700 7.670 1.180 ;
        RECT  9.670 0.300 9.870 1.180 ;
        RECT  10.160 0.300 12.290 0.460 ;
        RECT  12.110 0.300 12.290 0.960 ;
        RECT  12.110 0.800 12.830 0.960 ;
        RECT  12.670 0.800 12.830 1.270 ;
        RECT  10.160 0.300 10.430 1.780 ;
        RECT  13.060 0.400 13.320 1.600 ;
        RECT  13.060 0.950 14.220 1.230 ;
        RECT  12.110 1.120 12.390 1.600 ;
        RECT  13.060 0.950 13.330 1.600 ;
        RECT  12.110 1.440 13.330 1.600 ;
        RECT  14.900 1.050 15.760 1.280 ;
        RECT  10.860 1.330 11.950 1.610 ;
        RECT  11.670 0.620 11.950 1.920 ;
        RECT  14.900 1.050 15.080 1.920 ;
        RECT  11.560 1.760 15.080 1.920 ;
        RECT  11.560 1.330 11.860 2.100 ;
        LAYER VTPH ;
        RECT  6.250 0.970 7.370 2.400 ;
        RECT  0.420 1.040 1.750 2.400 ;
        RECT  10.180 1.020 11.400 2.400 ;
        RECT  9.730 1.090 11.400 2.400 ;
        RECT  12.860 1.080 14.680 2.400 ;
        RECT  6.250 1.060 8.070 2.400 ;
        RECT  0.000 1.140 8.070 2.400 ;
        RECT  9.730 1.140 16.400 2.400 ;
        RECT  0.000 1.180 16.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.400 0.970 ;
        RECT  7.370 0.000 16.400 1.020 ;
        RECT  0.000 0.000 6.250 1.040 ;
        RECT  7.370 0.000 10.180 1.060 ;
        RECT  11.400 0.000 16.400 1.080 ;
        RECT  8.070 0.000 10.180 1.090 ;
        RECT  0.000 0.000 0.420 1.140 ;
        RECT  1.750 0.000 6.250 1.140 ;
        RECT  11.400 0.000 12.860 1.140 ;
        RECT  14.680 0.000 16.400 1.140 ;
        RECT  8.070 0.000 9.730 1.180 ;
    END
END DFEZRM4HM

MACRO DFEZRM2HM
    CLASS CORE ;
    FOREIGN DFEZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        ANTENNAGATEAREA 0.089  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.036  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.950 1.900 1.150 ;
        LAYER ME2 ;
        RECT  1.700 0.700 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.500 0.950 2.080 1.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        ANTENNAGATEAREA 0.059  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.898  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.180 1.050 4.380 1.250 ;
        LAYER ME2 ;
        RECT  4.100 0.810 4.380 1.610 ;
        LAYER ME1 ;
        RECT  4.180 0.940 4.540 1.360 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.530 1.400 13.960 1.600 ;
        RECT  13.780 0.400 13.960 1.600 ;
        RECT  13.630 0.400 13.960 0.770 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.690 1.440 15.100 2.100 ;
        RECT  14.900 0.400 15.100 2.100 ;
        RECT  14.690 0.400 15.100 0.710 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        ANTENNAGATEAREA 0.220  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.729  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 0.950 0.700 1.150 ;
        LAYER ME2 ;
        RECT  0.500 0.700 0.700 1.340 ;
        LAYER ME1 ;
        RECT  0.500 0.810 0.760 1.280 ;
        END
    END E
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.110  LAYER ME1  ;
        ANTENNAGATEAREA 0.110  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.486  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.220 1.260 3.420 1.460 ;
        LAYER ME2 ;
        RECT  3.220 0.810 3.500 1.610 ;
        LAYER ME1 ;
        RECT  3.120 1.260 3.520 1.600 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.130 2.080 14.410 2.540 ;
        RECT  12.450 2.080 12.730 2.540 ;
        RECT  7.930 1.860 8.210 2.540 ;
        RECT  4.070 1.860 4.350 2.540 ;
        RECT  2.680 2.080 2.960 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.230 -0.140 14.430 0.720 ;
        RECT  12.550 -0.140 12.710 0.600 ;
        RECT  8.390 -0.140 8.670 0.540 ;
        RECT  3.580 -0.140 3.800 0.410 ;
        RECT  0.620 -0.140 0.900 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.960 0.910 1.160 1.600 ;
        RECT  2.260 0.940 2.460 1.600 ;
        RECT  0.140 1.440 2.460 1.600 ;
        RECT  0.140 0.410 0.340 2.030 ;
        RECT  1.100 0.300 3.310 0.460 ;
        RECT  1.100 0.300 1.380 0.590 ;
        RECT  2.760 0.940 3.990 1.100 ;
        RECT  3.770 0.940 3.990 1.340 ;
        RECT  2.760 0.940 2.960 1.500 ;
        RECT  4.770 0.620 5.060 0.840 ;
        RECT  4.830 0.620 5.060 1.250 ;
        RECT  4.830 0.970 5.570 1.250 ;
        RECT  4.830 0.620 5.030 1.760 ;
        RECT  5.690 0.620 5.970 0.820 ;
        RECT  5.770 0.930 6.070 1.220 ;
        RECT  5.770 0.620 5.970 1.730 ;
        RECT  3.960 0.300 6.410 0.460 ;
        RECT  6.210 0.300 6.410 0.600 ;
        RECT  3.960 0.300 4.120 0.780 ;
        RECT  1.880 0.620 4.120 0.780 ;
        RECT  3.750 1.540 4.670 1.700 ;
        RECT  3.750 1.540 3.910 1.920 ;
        RECT  1.660 1.760 3.910 1.920 ;
        RECT  4.510 1.540 4.670 2.100 ;
        RECT  1.660 1.760 1.860 2.080 ;
        RECT  6.320 1.480 6.520 2.100 ;
        RECT  4.510 1.940 6.520 2.100 ;
        RECT  6.880 0.370 7.190 0.710 ;
        RECT  6.880 0.370 7.080 1.650 ;
        RECT  6.880 1.490 8.710 1.650 ;
        RECT  8.490 1.490 8.710 1.840 ;
        RECT  9.180 0.660 9.460 1.180 ;
        RECT  8.090 1.020 9.460 1.180 ;
        RECT  9.300 0.660 9.460 1.760 ;
        RECT  9.300 1.480 9.530 1.760 ;
        RECT  8.850 0.300 9.870 0.460 ;
        RECT  8.850 0.300 9.020 0.860 ;
        RECT  7.470 0.700 9.020 0.860 ;
        RECT  7.470 0.700 7.670 1.180 ;
        RECT  9.670 0.300 9.870 1.180 ;
        RECT  10.160 0.300 12.290 0.460 ;
        RECT  12.110 0.300 12.290 0.960 ;
        RECT  12.110 0.800 12.830 0.960 ;
        RECT  12.670 0.800 12.830 1.270 ;
        RECT  10.160 0.300 10.430 1.780 ;
        RECT  13.060 0.400 13.320 1.600 ;
        RECT  13.060 0.950 13.470 1.230 ;
        RECT  12.110 1.120 12.390 1.600 ;
        RECT  13.060 0.950 13.330 1.600 ;
        RECT  12.110 1.440 13.330 1.600 ;
        RECT  14.220 0.980 14.540 1.280 ;
        RECT  10.860 1.330 11.950 1.610 ;
        RECT  11.670 0.620 11.950 1.920 ;
        RECT  14.220 0.980 14.400 1.920 ;
        RECT  11.560 1.760 14.400 1.920 ;
        RECT  11.560 1.330 11.860 2.100 ;
        LAYER VTPH ;
        RECT  6.250 0.970 7.370 2.400 ;
        RECT  0.420 1.040 1.750 2.400 ;
        RECT  10.180 1.020 11.400 2.400 ;
        RECT  9.730 1.090 11.400 2.400 ;
        RECT  12.860 1.080 14.040 2.400 ;
        RECT  6.250 1.060 8.070 2.400 ;
        RECT  0.000 1.140 8.070 2.400 ;
        RECT  9.730 1.140 15.200 2.400 ;
        RECT  0.000 1.180 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 0.970 ;
        RECT  7.370 0.000 15.200 1.020 ;
        RECT  0.000 0.000 6.250 1.040 ;
        RECT  7.370 0.000 10.180 1.060 ;
        RECT  11.400 0.000 15.200 1.080 ;
        RECT  8.070 0.000 10.180 1.090 ;
        RECT  0.000 0.000 0.420 1.140 ;
        RECT  1.750 0.000 6.250 1.140 ;
        RECT  11.400 0.000 12.860 1.140 ;
        RECT  14.040 0.000 15.200 1.140 ;
        RECT  8.070 0.000 9.730 1.180 ;
    END
END DFEZRM2HM

MACRO DFEZRM1HM
    CLASS CORE ;
    FOREIGN DFEZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.823  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 0.950 1.900 1.150 ;
        LAYER ME2 ;
        RECT  1.700 0.700 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.500 0.950 2.080 1.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.049  LAYER ME1  ;
        ANTENNAGATEAREA 0.049  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.244  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.180 1.050 4.380 1.250 ;
        LAYER ME2 ;
        RECT  4.100 0.810 4.380 1.610 ;
        LAYER ME1 ;
        RECT  4.180 0.940 4.540 1.360 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.332  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.530 1.400 13.960 1.600 ;
        RECT  13.790 0.360 13.960 1.600 ;
        RECT  13.630 0.360 13.960 0.770 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.690 1.550 15.100 1.830 ;
        RECT  14.900 0.390 15.100 1.830 ;
        RECT  14.690 0.390 15.100 0.670 ;
        END
    END QB
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        ANTENNAGATEAREA 0.161  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.361  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 0.950 0.700 1.150 ;
        LAYER ME2 ;
        RECT  0.500 0.700 0.700 1.340 ;
        LAYER ME1 ;
        RECT  0.500 0.810 0.760 1.280 ;
        END
    END E
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.010  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.220 1.260 3.420 1.460 ;
        LAYER ME2 ;
        RECT  3.220 0.810 3.500 1.610 ;
        LAYER ME1 ;
        RECT  3.120 1.260 3.520 1.600 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.130 2.080 14.410 2.540 ;
        RECT  12.450 2.080 12.730 2.540 ;
        RECT  7.930 1.860 8.210 2.540 ;
        RECT  4.070 1.860 4.350 2.540 ;
        RECT  2.680 2.080 2.960 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.230 -0.140 14.430 0.650 ;
        RECT  12.550 -0.140 12.710 0.640 ;
        RECT  8.390 -0.140 8.670 0.540 ;
        RECT  3.580 -0.140 3.800 0.410 ;
        RECT  0.620 -0.140 0.900 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.960 0.910 1.160 1.600 ;
        RECT  2.260 0.940 2.460 1.600 ;
        RECT  0.140 1.440 2.460 1.600 ;
        RECT  0.140 0.340 0.340 2.030 ;
        RECT  1.100 0.300 3.310 0.460 ;
        RECT  1.100 0.300 1.380 0.590 ;
        RECT  2.760 0.940 3.990 1.100 ;
        RECT  3.770 0.940 3.990 1.340 ;
        RECT  2.760 0.940 2.960 1.500 ;
        RECT  4.770 0.620 5.060 0.840 ;
        RECT  4.830 0.620 5.060 1.250 ;
        RECT  4.830 0.970 5.570 1.250 ;
        RECT  4.830 0.620 5.030 1.760 ;
        RECT  5.690 0.620 5.970 0.820 ;
        RECT  5.770 0.930 6.070 1.220 ;
        RECT  5.770 0.620 5.970 1.730 ;
        RECT  3.960 0.300 6.410 0.460 ;
        RECT  6.210 0.300 6.410 0.600 ;
        RECT  3.960 0.300 4.120 0.780 ;
        RECT  1.880 0.620 4.120 0.780 ;
        RECT  3.750 1.540 4.670 1.700 ;
        RECT  3.750 1.540 3.910 1.920 ;
        RECT  1.660 1.760 3.910 1.920 ;
        RECT  4.510 1.540 4.670 2.100 ;
        RECT  1.660 1.760 1.860 2.080 ;
        RECT  6.320 1.480 6.520 2.100 ;
        RECT  4.510 1.940 6.520 2.100 ;
        RECT  6.860 0.390 7.140 1.650 ;
        RECT  6.860 1.490 8.710 1.650 ;
        RECT  8.490 1.490 8.710 1.840 ;
        RECT  9.180 0.660 9.460 1.180 ;
        RECT  8.090 1.020 9.460 1.180 ;
        RECT  9.300 0.660 9.460 1.760 ;
        RECT  9.300 1.480 9.530 1.760 ;
        RECT  8.850 0.300 9.870 0.460 ;
        RECT  8.850 0.300 9.020 0.860 ;
        RECT  7.470 0.700 9.020 0.860 ;
        RECT  7.470 0.700 7.670 1.180 ;
        RECT  9.670 0.300 9.870 1.180 ;
        RECT  10.160 0.300 12.290 0.460 ;
        RECT  12.110 0.300 12.290 0.960 ;
        RECT  12.110 0.800 12.830 0.960 ;
        RECT  12.670 0.800 12.830 1.270 ;
        RECT  10.160 0.300 10.430 1.780 ;
        RECT  13.060 0.370 13.320 1.600 ;
        RECT  13.060 0.950 13.470 1.230 ;
        RECT  12.110 1.120 12.390 1.600 ;
        RECT  13.060 0.950 13.330 1.600 ;
        RECT  12.110 1.440 13.330 1.600 ;
        RECT  14.220 0.980 14.540 1.280 ;
        RECT  10.860 1.330 11.950 1.610 ;
        RECT  11.670 0.620 11.950 1.920 ;
        RECT  14.220 0.980 14.400 1.920 ;
        RECT  11.560 1.760 14.400 1.920 ;
        RECT  11.560 1.330 11.840 2.100 ;
        LAYER VTPH ;
        RECT  6.270 0.910 7.320 2.400 ;
        RECT  6.270 0.990 7.370 2.400 ;
        RECT  0.420 1.040 1.750 2.400 ;
        RECT  6.230 1.100 8.070 2.400 ;
        RECT  10.180 1.020 11.400 2.400 ;
        RECT  9.730 1.090 11.400 2.400 ;
        RECT  12.860 1.080 14.040 2.400 ;
        RECT  6.270 1.060 8.070 2.400 ;
        RECT  0.000 1.140 8.070 2.400 ;
        RECT  9.730 1.140 15.200 2.400 ;
        RECT  0.000 1.180 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 0.910 ;
        RECT  7.320 0.000 15.200 0.990 ;
        RECT  7.370 0.000 15.200 1.020 ;
        RECT  0.000 0.000 6.270 1.040 ;
        RECT  7.370 0.000 10.180 1.060 ;
        RECT  11.400 0.000 15.200 1.080 ;
        RECT  8.070 0.000 10.180 1.090 ;
        RECT  1.750 0.000 6.270 1.100 ;
        RECT  0.000 0.000 0.420 1.140 ;
        RECT  1.750 0.000 6.230 1.140 ;
        RECT  11.400 0.000 12.860 1.140 ;
        RECT  14.040 0.000 15.200 1.140 ;
        RECT  8.070 0.000 9.730 1.180 ;
    END
END DFEZRM1HM

MACRO DFERM8HM
    CLASS CORE ;
    FOREIGN DFERM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        ANTENNAGATEAREA 0.120  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.110 3.500 1.310 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.620 1.080 3.820 1.460 ;
        RECT  3.200 1.080 3.820 1.340 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.097  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.100 1.360 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.840 0.700 1.360 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.968  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.180 1.400 17.660 1.600 ;
        RECT  17.300 0.420 17.660 1.600 ;
        RECT  16.380 1.230 17.660 1.600 ;
        RECT  16.380 0.420 16.540 1.600 ;
        RECT  16.180 0.420 16.540 0.700 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.986  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  19.500 0.440 19.700 2.100 ;
        RECT  18.460 0.900 19.700 1.170 ;
        RECT  18.460 0.440 18.730 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.650 1.120 15.680 1.280 ;
        RECT  15.460 1.000 15.680 1.280 ;
        RECT  12.840 0.980 13.940 1.140 ;
        RECT  11.700 1.400 13.000 1.560 ;
        RECT  12.840 0.980 13.000 1.560 ;
        RECT  9.650 1.940 11.900 2.100 ;
        RECT  11.700 1.400 11.900 2.100 ;
        RECT  9.650 1.540 9.810 2.100 ;
        RECT  8.890 1.540 9.810 1.700 ;
        RECT  8.890 1.540 9.050 2.020 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 20.400 2.540 ;
        RECT  20.020 1.480 20.220 2.540 ;
        RECT  18.980 1.460 19.180 2.540 ;
        RECT  17.860 2.080 18.140 2.540 ;
        RECT  16.740 2.080 17.020 2.540 ;
        RECT  15.600 2.080 15.880 2.540 ;
        RECT  13.280 2.080 13.560 2.540 ;
        RECT  9.210 1.860 9.490 2.540 ;
        RECT  7.550 1.860 7.830 2.540 ;
        RECT  2.920 1.820 3.120 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 20.400 0.140 ;
        RECT  20.020 -0.140 20.220 0.720 ;
        RECT  18.980 -0.140 19.180 0.720 ;
        RECT  17.860 -0.140 18.140 0.700 ;
        RECT  16.740 -0.140 17.020 0.650 ;
        RECT  15.640 -0.140 15.920 0.500 ;
        RECT  13.440 -0.140 13.720 0.320 ;
        RECT  9.070 -0.140 9.350 0.550 ;
        RECT  3.240 -0.140 3.500 0.600 ;
        RECT  0.700 -0.140 0.980 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.360 2.060 0.560 ;
        RECT  1.420 0.360 1.580 1.750 ;
        RECT  0.100 0.300 0.380 0.580 ;
        RECT  1.740 0.890 2.760 1.190 ;
        RECT  0.100 0.300 0.270 2.080 ;
        RECT  0.100 1.520 1.260 1.680 ;
        RECT  1.100 1.520 1.260 2.100 ;
        RECT  0.100 1.520 0.380 2.080 ;
        RECT  1.740 0.890 1.900 2.100 ;
        RECT  1.100 1.940 1.900 2.100 ;
        RECT  3.980 0.680 4.920 0.950 ;
        RECT  4.700 0.680 4.920 1.340 ;
        RECT  3.980 0.680 4.140 1.780 ;
        RECT  3.710 1.620 4.140 1.780 ;
        RECT  5.080 0.670 5.360 1.780 ;
        RECT  5.080 1.350 5.520 1.780 ;
        RECT  4.880 1.560 5.520 1.780 ;
        RECT  3.660 0.300 5.840 0.460 ;
        RECT  2.300 0.380 3.080 0.600 ;
        RECT  5.560 0.300 5.840 0.710 ;
        RECT  2.920 0.380 3.080 0.920 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  2.920 0.760 3.820 0.920 ;
        RECT  2.060 1.500 3.460 1.660 ;
        RECT  3.300 1.500 3.460 2.100 ;
        RECT  2.060 1.500 2.220 2.100 ;
        RECT  5.680 1.640 5.970 2.100 ;
        RECT  3.300 1.940 5.970 2.100 ;
        RECT  6.210 0.410 6.440 0.740 ;
        RECT  6.210 0.550 7.010 0.740 ;
        RECT  6.850 0.550 7.010 1.020 ;
        RECT  8.150 0.770 8.430 1.020 ;
        RECT  6.850 0.860 8.430 1.020 ;
        RECT  6.210 0.410 6.370 1.940 ;
        RECT  6.210 1.740 6.610 1.940 ;
        RECT  6.930 1.540 8.730 1.700 ;
        RECT  8.450 1.540 8.730 1.860 ;
        RECT  6.930 1.540 7.230 1.970 ;
        RECT  6.530 0.900 6.690 1.380 ;
        RECT  10.100 1.030 10.380 1.380 ;
        RECT  6.530 1.220 10.380 1.380 ;
        RECT  7.170 0.420 8.800 0.580 ;
        RECT  7.170 0.420 7.450 0.640 ;
        RECT  9.770 0.500 10.060 0.870 ;
        RECT  9.770 0.710 10.700 0.870 ;
        RECT  8.640 0.420 8.800 1.060 ;
        RECT  9.770 0.500 9.930 1.060 ;
        RECT  8.640 0.900 9.930 1.060 ;
        RECT  10.540 0.710 10.700 1.780 ;
        RECT  9.970 1.620 10.700 1.780 ;
        RECT  11.240 0.860 11.460 1.200 ;
        RECT  11.240 1.040 12.310 1.200 ;
        RECT  12.680 0.620 12.960 0.820 ;
        RECT  11.800 0.660 12.960 0.820 ;
        RECT  12.480 0.660 12.680 1.220 ;
        RECT  10.860 0.300 13.280 0.460 ;
        RECT  13.120 0.300 13.280 0.660 ;
        RECT  13.120 0.500 14.350 0.660 ;
        RECT  14.190 0.500 14.350 0.920 ;
        RECT  14.190 0.720 14.840 0.920 ;
        RECT  10.860 0.300 11.020 1.780 ;
        RECT  10.860 1.580 11.220 1.780 ;
        RECT  14.710 0.340 15.170 0.520 ;
        RECT  15.010 0.340 15.170 0.840 ;
        RECT  15.010 0.680 16.020 0.840 ;
        RECT  15.860 0.960 16.220 1.240 ;
        RECT  13.160 1.320 13.440 1.600 ;
        RECT  15.860 0.680 16.020 1.600 ;
        RECT  13.160 1.440 16.020 1.600 ;
        RECT  12.300 1.720 12.580 1.920 ;
        RECT  18.050 1.050 18.270 1.920 ;
        RECT  12.300 1.760 18.270 1.920 ;
        LAYER VTPH ;
        RECT  0.400 1.000 2.250 2.400 ;
        RECT  13.200 1.080 18.220 2.400 ;
        RECT  0.400 1.100 2.930 2.400 ;
        RECT  0.000 1.140 2.930 2.400 ;
        RECT  8.330 1.110 10.210 2.400 ;
        RECT  12.430 1.140 20.400 2.400 ;
        RECT  0.000 1.260 20.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 20.400 1.000 ;
        RECT  2.250 0.000 20.400 1.080 ;
        RECT  2.250 0.000 13.200 1.100 ;
        RECT  2.930 0.000 13.200 1.110 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  10.210 0.000 13.200 1.140 ;
        RECT  18.220 0.000 20.400 1.140 ;
        RECT  2.930 0.000 8.330 1.260 ;
        RECT  10.210 0.000 12.430 1.260 ;
    END
END DFERM8HM

MACRO DFERM4HM
    CLASS CORE ;
    FOREIGN DFERM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        ANTENNAGATEAREA 0.060  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.110 3.500 1.310 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.620 1.080 3.820 1.460 ;
        RECT  3.200 1.080 3.820 1.340 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.100 1.360 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.840 0.700 1.360 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.980 1.400 16.380 1.600 ;
        RECT  16.180 0.420 16.380 1.600 ;
        RECT  15.980 0.420 16.380 0.700 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.490  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.140 0.440 17.500 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.450 1.120 15.480 1.280 ;
        RECT  15.260 1.000 15.480 1.280 ;
        RECT  12.650 0.980 13.740 1.140 ;
        RECT  11.300 1.400 12.810 1.560 ;
        RECT  12.650 0.980 12.810 1.560 ;
        RECT  9.470 1.940 11.500 2.100 ;
        RECT  11.300 1.400 11.500 2.100 ;
        RECT  9.470 1.540 9.630 2.100 ;
        RECT  8.710 1.540 9.630 1.700 ;
        RECT  8.710 1.540 8.870 2.020 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.000 2.540 ;
        RECT  17.660 1.470 17.860 2.540 ;
        RECT  16.540 2.080 16.820 2.540 ;
        RECT  15.400 2.080 15.680 2.540 ;
        RECT  13.100 2.080 13.380 2.540 ;
        RECT  9.030 1.860 9.310 2.540 ;
        RECT  7.370 1.860 7.650 2.540 ;
        RECT  2.920 1.820 3.120 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.000 0.140 ;
        RECT  17.660 -0.140 17.860 0.720 ;
        RECT  16.540 -0.140 16.820 0.500 ;
        RECT  15.440 -0.140 15.720 0.500 ;
        RECT  13.260 -0.140 13.480 0.380 ;
        RECT  8.890 -0.140 9.170 0.550 ;
        RECT  3.240 -0.140 3.500 0.600 ;
        RECT  0.700 -0.140 0.980 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.360 2.060 0.560 ;
        RECT  1.420 0.360 1.580 1.750 ;
        RECT  0.100 0.300 0.380 0.580 ;
        RECT  1.740 0.860 2.760 1.140 ;
        RECT  0.100 0.300 0.270 2.080 ;
        RECT  0.100 1.520 1.260 1.680 ;
        RECT  1.100 1.520 1.260 2.100 ;
        RECT  0.100 1.520 0.380 2.080 ;
        RECT  1.740 0.860 1.900 2.100 ;
        RECT  1.100 1.940 1.900 2.100 ;
        RECT  3.980 0.650 4.200 1.340 ;
        RECT  3.980 1.060 4.740 1.340 ;
        RECT  3.980 0.650 4.140 1.780 ;
        RECT  3.710 1.620 4.140 1.780 ;
        RECT  4.900 0.700 5.180 1.780 ;
        RECT  4.900 1.350 5.340 1.780 ;
        RECT  4.700 1.560 5.340 1.780 ;
        RECT  3.660 0.300 5.660 0.460 ;
        RECT  2.300 0.380 3.080 0.600 ;
        RECT  5.380 0.300 5.660 0.710 ;
        RECT  2.920 0.380 3.080 0.920 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  2.920 0.760 3.820 0.920 ;
        RECT  2.060 1.500 3.460 1.660 ;
        RECT  3.300 1.500 3.460 2.100 ;
        RECT  2.060 1.500 2.220 2.100 ;
        RECT  5.500 1.640 5.790 2.100 ;
        RECT  3.300 1.940 5.790 2.100 ;
        RECT  6.030 0.410 6.830 0.740 ;
        RECT  6.670 0.410 6.830 1.020 ;
        RECT  7.970 0.770 8.250 1.020 ;
        RECT  6.670 0.860 8.250 1.020 ;
        RECT  6.030 0.410 6.190 1.940 ;
        RECT  6.030 1.740 6.430 1.940 ;
        RECT  6.750 1.540 8.550 1.700 ;
        RECT  8.270 1.540 8.550 1.860 ;
        RECT  6.750 1.540 7.050 1.970 ;
        RECT  6.350 0.900 6.510 1.380 ;
        RECT  9.890 1.030 10.170 1.380 ;
        RECT  6.350 1.220 10.170 1.380 ;
        RECT  6.990 0.420 8.620 0.580 ;
        RECT  6.990 0.420 7.270 0.640 ;
        RECT  9.660 0.500 9.940 0.870 ;
        RECT  9.390 0.700 9.940 0.870 ;
        RECT  9.390 0.710 10.490 0.870 ;
        RECT  8.460 0.420 8.620 1.060 ;
        RECT  9.390 0.700 9.550 1.060 ;
        RECT  8.460 0.900 9.550 1.060 ;
        RECT  10.330 0.710 10.490 1.780 ;
        RECT  9.790 1.620 10.490 1.780 ;
        RECT  11.050 0.860 11.270 1.200 ;
        RECT  11.050 1.040 12.120 1.200 ;
        RECT  12.490 0.620 12.770 0.820 ;
        RECT  11.610 0.660 12.770 0.820 ;
        RECT  12.290 0.660 12.490 1.220 ;
        RECT  10.670 0.300 13.090 0.460 ;
        RECT  12.930 0.300 13.090 0.820 ;
        RECT  12.930 0.660 14.150 0.820 ;
        RECT  13.990 0.720 14.640 0.920 ;
        RECT  10.670 0.300 10.830 1.780 ;
        RECT  10.670 1.580 11.030 1.780 ;
        RECT  14.510 0.340 14.970 0.520 ;
        RECT  14.810 0.340 14.970 0.840 ;
        RECT  14.810 0.680 15.820 0.840 ;
        RECT  15.660 0.960 16.020 1.240 ;
        RECT  12.970 1.320 13.250 1.600 ;
        RECT  15.660 0.680 15.820 1.600 ;
        RECT  12.970 1.440 15.820 1.600 ;
        RECT  12.110 1.720 12.390 1.920 ;
        RECT  16.730 1.050 16.950 1.920 ;
        RECT  12.110 1.760 16.950 1.920 ;
        LAYER VTPH ;
        RECT  0.400 1.000 2.250 2.400 ;
        RECT  13.010 1.080 16.900 2.400 ;
        RECT  0.400 1.100 2.930 2.400 ;
        RECT  0.000 1.140 2.930 2.400 ;
        RECT  8.150 1.110 10.030 2.400 ;
        RECT  12.240 1.140 18.000 2.400 ;
        RECT  0.000 1.260 18.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.000 1.000 ;
        RECT  2.250 0.000 18.000 1.080 ;
        RECT  2.250 0.000 13.010 1.100 ;
        RECT  2.930 0.000 13.010 1.110 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  10.030 0.000 13.010 1.140 ;
        RECT  16.900 0.000 18.000 1.140 ;
        RECT  2.930 0.000 8.150 1.260 ;
        RECT  10.030 0.000 12.240 1.260 ;
    END
END DFERM4HM

MACRO DFERM2HM
    CLASS CORE ;
    FOREIGN DFERM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.060  LAYER ME1  ;
        ANTENNAGATEAREA 0.060  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.667  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.110 3.500 1.310 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.620 1.080 3.820 1.460 ;
        RECT  3.200 1.080 3.820 1.340 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.100 1.360 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.840 0.700 1.360 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.448  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.780 0.420 15.160 0.760 ;
        RECT  14.740 1.400 15.020 1.600 ;
        RECT  14.780 0.420 15.020 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.000 0.440 16.300 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.420 0.820 13.650 1.280 ;
        RECT  12.680 0.820 13.650 0.980 ;
        RECT  11.300 1.400 12.840 1.560 ;
        RECT  12.680 0.820 12.840 1.560 ;
        RECT  9.550 1.940 11.500 2.100 ;
        RECT  11.300 1.400 11.500 2.100 ;
        RECT  9.550 1.540 9.710 2.100 ;
        RECT  8.730 1.540 9.710 1.700 ;
        RECT  8.730 1.400 9.010 1.700 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.400 2.540 ;
        RECT  15.500 1.460 15.700 2.540 ;
        RECT  14.210 2.080 14.490 2.540 ;
        RECT  12.920 2.080 13.200 2.540 ;
        RECT  8.990 1.860 9.270 2.540 ;
        RECT  7.370 1.860 7.650 2.540 ;
        RECT  2.920 1.820 3.120 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.400 0.140 ;
        RECT  15.460 -0.140 15.680 0.700 ;
        RECT  13.000 -0.140 13.280 0.320 ;
        RECT  8.800 -0.140 9.080 0.540 ;
        RECT  3.240 -0.140 3.500 0.600 ;
        RECT  0.700 -0.140 0.980 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.360 2.060 0.560 ;
        RECT  1.420 0.360 1.580 1.750 ;
        RECT  0.100 0.300 0.380 0.580 ;
        RECT  1.740 0.860 2.760 1.140 ;
        RECT  0.100 0.300 0.270 2.080 ;
        RECT  0.100 1.520 1.260 1.680 ;
        RECT  1.100 1.520 1.260 2.100 ;
        RECT  0.100 1.520 0.380 2.080 ;
        RECT  1.740 0.860 1.900 2.100 ;
        RECT  1.100 1.940 1.900 2.100 ;
        RECT  3.980 0.650 4.200 1.340 ;
        RECT  3.980 1.060 4.740 1.340 ;
        RECT  3.980 0.650 4.140 1.780 ;
        RECT  3.710 1.620 4.140 1.780 ;
        RECT  4.900 0.700 5.180 1.780 ;
        RECT  4.900 1.460 5.340 1.780 ;
        RECT  4.700 1.560 5.340 1.780 ;
        RECT  3.660 0.300 5.660 0.460 ;
        RECT  2.300 0.380 3.080 0.600 ;
        RECT  5.380 0.300 5.660 0.710 ;
        RECT  2.920 0.380 3.080 0.920 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  2.920 0.760 3.820 0.920 ;
        RECT  2.060 1.500 3.460 1.660 ;
        RECT  3.300 1.500 3.460 2.100 ;
        RECT  2.060 1.500 2.220 2.100 ;
        RECT  5.500 1.640 5.790 2.100 ;
        RECT  3.300 1.940 5.790 2.100 ;
        RECT  6.750 1.540 8.130 1.700 ;
        RECT  7.850 1.540 8.130 1.860 ;
        RECT  6.750 1.540 7.050 1.910 ;
        RECT  6.030 0.410 6.830 0.740 ;
        RECT  6.670 0.410 6.830 1.020 ;
        RECT  7.950 0.770 8.230 1.020 ;
        RECT  6.670 0.860 8.230 1.020 ;
        RECT  6.030 0.410 6.190 1.940 ;
        RECT  6.030 1.740 6.430 1.940 ;
        RECT  6.350 0.900 6.510 1.380 ;
        RECT  8.390 1.020 9.910 1.220 ;
        RECT  9.690 1.020 9.910 1.310 ;
        RECT  6.350 1.220 8.550 1.380 ;
        RECT  6.990 0.420 8.550 0.580 ;
        RECT  6.990 0.420 7.270 0.640 ;
        RECT  8.390 0.420 8.550 0.860 ;
        RECT  9.410 0.500 9.690 0.860 ;
        RECT  8.390 0.700 10.260 0.860 ;
        RECT  10.100 0.700 10.260 1.780 ;
        RECT  9.880 1.580 10.260 1.780 ;
        RECT  10.800 0.860 11.020 1.200 ;
        RECT  10.800 1.040 11.870 1.200 ;
        RECT  11.440 0.620 12.520 0.820 ;
        RECT  12.040 0.620 12.240 1.220 ;
        RECT  10.420 0.300 12.840 0.460 ;
        RECT  12.680 0.300 12.840 0.660 ;
        RECT  12.680 0.500 13.970 0.660 ;
        RECT  13.810 0.500 13.970 1.280 ;
        RECT  13.810 0.960 14.130 1.280 ;
        RECT  10.420 0.300 10.580 1.780 ;
        RECT  10.420 1.580 10.780 1.780 ;
        RECT  14.180 0.340 14.450 0.700 ;
        RECT  14.290 0.960 14.610 1.240 ;
        RECT  13.000 1.140 13.220 1.600 ;
        RECT  14.290 0.340 14.450 1.600 ;
        RECT  13.000 1.440 14.450 1.600 ;
        RECT  15.180 0.940 15.720 1.220 ;
        RECT  11.860 1.720 12.140 1.920 ;
        RECT  15.180 0.940 15.340 1.920 ;
        RECT  11.860 1.760 15.340 1.920 ;
        LAYER VTPH ;
        RECT  0.400 1.000 2.250 2.400 ;
        RECT  12.760 1.080 15.680 2.400 ;
        RECT  0.400 1.100 2.930 2.400 ;
        RECT  0.000 1.140 2.930 2.400 ;
        RECT  8.130 1.110 10.400 2.400 ;
        RECT  11.990 1.140 16.400 2.400 ;
        RECT  0.000 1.260 16.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.400 1.000 ;
        RECT  2.250 0.000 16.400 1.080 ;
        RECT  2.250 0.000 12.760 1.100 ;
        RECT  2.930 0.000 12.760 1.110 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  10.400 0.000 12.760 1.140 ;
        RECT  15.680 0.000 16.400 1.140 ;
        RECT  2.930 0.000 8.130 1.260 ;
        RECT  10.400 0.000 11.990 1.260 ;
    END
END DFERM2HM

MACRO DFERM1HM
    CLASS CORE ;
    FOREIGN DFERM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.058  LAYER ME1  ;
        ANTENNAGATEAREA 0.058  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.028  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.110 3.500 1.310 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.620 1.080 3.820 1.460 ;
        RECT  3.200 1.080 3.820 1.340 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.100 1.360 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.148  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.460 0.840 0.700 1.360 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.331  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.780 0.420 15.160 0.760 ;
        RECT  14.740 1.400 15.020 1.600 ;
        RECT  14.780 0.420 15.020 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  16.000 0.440 16.300 2.100 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.420 0.820 13.650 1.280 ;
        RECT  12.680 0.820 13.650 0.980 ;
        RECT  11.300 1.400 12.840 1.560 ;
        RECT  12.680 0.820 12.840 1.560 ;
        RECT  9.550 1.940 11.500 2.100 ;
        RECT  11.300 1.400 11.500 2.100 ;
        RECT  9.550 1.540 9.710 2.100 ;
        RECT  8.730 1.540 9.710 1.700 ;
        RECT  8.730 1.400 9.010 1.700 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.400 2.540 ;
        RECT  15.500 1.460 15.700 2.540 ;
        RECT  14.210 2.080 14.490 2.540 ;
        RECT  12.920 2.080 13.200 2.540 ;
        RECT  8.990 1.860 9.270 2.540 ;
        RECT  7.370 1.860 7.650 2.540 ;
        RECT  2.920 1.820 3.120 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.400 0.140 ;
        RECT  15.460 -0.140 15.680 0.700 ;
        RECT  13.000 -0.140 13.280 0.320 ;
        RECT  8.800 -0.140 9.080 0.540 ;
        RECT  3.240 -0.140 3.500 0.600 ;
        RECT  0.700 -0.140 0.980 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.420 0.360 2.060 0.560 ;
        RECT  1.420 0.360 1.580 1.660 ;
        RECT  0.100 0.340 0.380 0.620 ;
        RECT  1.740 0.860 2.760 1.140 ;
        RECT  0.100 0.340 0.270 2.080 ;
        RECT  0.100 1.520 1.260 1.680 ;
        RECT  1.100 1.520 1.260 2.100 ;
        RECT  0.100 1.520 0.380 2.080 ;
        RECT  1.740 0.860 1.900 2.100 ;
        RECT  1.100 1.940 1.900 2.100 ;
        RECT  3.980 0.650 4.200 1.340 ;
        RECT  3.980 1.060 4.740 1.340 ;
        RECT  3.980 0.650 4.140 1.780 ;
        RECT  3.710 1.620 4.140 1.780 ;
        RECT  4.900 0.700 5.180 1.780 ;
        RECT  4.900 1.460 5.340 1.780 ;
        RECT  4.700 1.560 5.340 1.780 ;
        RECT  3.660 0.300 5.660 0.460 ;
        RECT  2.300 0.380 3.080 0.580 ;
        RECT  5.380 0.300 5.660 0.710 ;
        RECT  2.920 0.380 3.080 0.920 ;
        RECT  3.660 0.300 3.820 0.920 ;
        RECT  2.920 0.760 3.820 0.920 ;
        RECT  2.060 1.500 3.460 1.660 ;
        RECT  2.060 1.500 2.220 1.890 ;
        RECT  3.300 1.500 3.460 2.100 ;
        RECT  5.500 1.640 5.790 2.100 ;
        RECT  3.300 1.940 5.790 2.100 ;
        RECT  6.750 1.540 8.130 1.700 ;
        RECT  7.850 1.540 8.130 1.860 ;
        RECT  6.750 1.540 7.050 1.910 ;
        RECT  6.030 0.410 6.830 0.740 ;
        RECT  6.670 0.410 6.830 1.020 ;
        RECT  7.950 0.770 8.230 1.020 ;
        RECT  6.670 0.860 8.230 1.020 ;
        RECT  6.030 0.410 6.190 1.940 ;
        RECT  6.030 1.740 6.430 1.940 ;
        RECT  6.350 0.900 6.510 1.380 ;
        RECT  8.390 1.020 9.910 1.220 ;
        RECT  9.690 1.020 9.910 1.310 ;
        RECT  6.350 1.220 8.550 1.380 ;
        RECT  6.990 0.420 8.550 0.580 ;
        RECT  6.990 0.420 7.270 0.640 ;
        RECT  8.390 0.420 8.550 0.860 ;
        RECT  9.410 0.500 9.690 0.860 ;
        RECT  8.390 0.700 10.260 0.860 ;
        RECT  10.100 0.700 10.260 1.780 ;
        RECT  9.880 1.580 10.260 1.780 ;
        RECT  10.800 0.860 11.020 1.200 ;
        RECT  10.800 1.040 11.870 1.200 ;
        RECT  11.440 0.620 12.520 0.820 ;
        RECT  12.040 0.620 12.240 1.220 ;
        RECT  10.420 0.300 12.840 0.460 ;
        RECT  12.680 0.300 12.840 0.660 ;
        RECT  12.680 0.500 13.970 0.660 ;
        RECT  13.810 0.500 13.970 1.280 ;
        RECT  13.810 0.960 14.130 1.280 ;
        RECT  10.420 0.300 10.580 1.780 ;
        RECT  10.420 1.580 10.780 1.780 ;
        RECT  14.180 0.340 14.450 0.670 ;
        RECT  14.290 0.960 14.610 1.240 ;
        RECT  13.000 1.140 13.220 1.600 ;
        RECT  14.290 0.340 14.450 1.600 ;
        RECT  13.000 1.440 14.450 1.600 ;
        RECT  15.180 0.940 15.720 1.220 ;
        RECT  11.860 1.720 12.140 1.920 ;
        RECT  15.180 0.940 15.340 1.920 ;
        RECT  11.860 1.760 15.340 1.920 ;
        LAYER VTPH ;
        RECT  0.400 1.000 2.250 2.400 ;
        RECT  12.760 1.080 15.680 2.400 ;
        RECT  0.400 1.100 2.930 2.400 ;
        RECT  0.000 1.140 2.930 2.400 ;
        RECT  8.130 1.110 10.400 2.400 ;
        RECT  11.990 1.140 16.400 2.400 ;
        RECT  0.000 1.260 16.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.400 1.000 ;
        RECT  2.250 0.000 16.400 1.080 ;
        RECT  2.250 0.000 12.760 1.100 ;
        RECT  2.930 0.000 12.760 1.110 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  10.400 0.000 12.760 1.140 ;
        RECT  15.680 0.000 16.400 1.140 ;
        RECT  2.930 0.000 8.130 1.260 ;
        RECT  10.400 0.000 11.990 1.260 ;
    END
END DFERM1HM

MACRO DFEQZRM8HM
    CLASS CORE ;
    FOREIGN DFEQZRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.054  LAYER ME1  ;
        ANTENNAGATEAREA 0.054  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.126  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 0.970 3.500 1.170 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.580 ;
        LAYER ME1 ;
        RECT  3.200 0.970 3.640 1.270 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 0.440 4.880 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.330 0.730 1.910 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.173  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.760 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.700 0.400 14.980 2.100 ;
        RECT  13.700 0.840 14.980 1.170 ;
        RECT  13.660 1.460 13.900 2.100 ;
        RECT  13.700 0.400 13.900 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  15.220 1.480 15.500 2.540 ;
        RECT  14.180 1.480 14.460 2.540 ;
        RECT  13.140 1.480 13.420 2.540 ;
        RECT  12.100 1.900 12.380 2.540 ;
        RECT  8.930 1.770 9.210 2.540 ;
        RECT  5.100 1.860 5.380 2.540 ;
        RECT  3.000 1.860 3.280 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  15.220 -0.140 15.500 0.680 ;
        RECT  14.180 -0.140 14.460 0.680 ;
        RECT  13.140 -0.140 13.420 0.670 ;
        RECT  12.160 -0.140 12.320 0.600 ;
        RECT  8.930 -0.140 9.210 0.320 ;
        RECT  5.580 -0.140 6.250 0.760 ;
        RECT  3.850 -0.140 4.130 0.320 ;
        RECT  0.620 -0.140 0.900 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.330 0.380 0.600 ;
        RECT  2.190 1.060 2.660 1.220 ;
        RECT  0.100 0.330 0.260 1.940 ;
        RECT  0.900 0.760 1.060 1.540 ;
        RECT  2.190 1.060 2.440 1.540 ;
        RECT  0.100 1.380 2.440 1.540 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.060 0.330 3.360 0.490 ;
        RECT  1.060 0.330 1.470 0.540 ;
        RECT  2.070 0.650 4.340 0.810 ;
        RECT  4.060 0.650 4.340 0.990 ;
        RECT  5.040 0.380 5.200 1.380 ;
        RECT  5.040 1.180 5.930 1.380 ;
        RECT  4.340 1.220 5.930 1.380 ;
        RECT  4.340 1.220 4.620 1.730 ;
        RECT  7.010 0.300 7.570 0.610 ;
        RECT  7.370 0.300 7.570 0.660 ;
        RECT  6.620 0.420 6.810 1.420 ;
        RECT  6.620 1.140 7.780 1.420 ;
        RECT  6.090 1.260 7.780 1.420 ;
        RECT  6.090 1.260 6.250 1.780 ;
        RECT  2.600 1.540 3.920 1.700 ;
        RECT  4.780 1.540 5.700 1.700 ;
        RECT  3.560 1.540 3.920 1.740 ;
        RECT  6.410 1.580 7.810 1.740 ;
        RECT  3.760 1.540 3.920 2.100 ;
        RECT  5.540 1.540 5.700 2.100 ;
        RECT  2.600 1.540 2.760 2.080 ;
        RECT  1.620 1.800 2.760 2.080 ;
        RECT  4.780 1.540 4.940 2.100 ;
        RECT  3.760 1.940 4.940 2.100 ;
        RECT  6.410 1.580 6.570 2.100 ;
        RECT  5.540 1.940 6.570 2.100 ;
        RECT  7.850 0.360 8.130 0.640 ;
        RECT  7.970 0.360 8.130 1.280 ;
        RECT  7.970 1.120 9.660 1.280 ;
        RECT  8.010 1.060 8.290 1.780 ;
        RECT  9.700 0.620 9.980 0.960 ;
        RECT  8.670 0.800 9.980 0.960 ;
        RECT  9.820 0.620 9.980 1.760 ;
        RECT  9.800 1.480 10.000 1.760 ;
        RECT  9.370 0.300 10.300 0.460 ;
        RECT  9.370 0.300 9.540 0.640 ;
        RECT  8.290 0.480 9.540 0.640 ;
        RECT  8.290 0.480 8.450 0.900 ;
        RECT  10.140 0.300 10.300 1.100 ;
        RECT  11.150 0.620 11.430 0.960 ;
        RECT  10.940 0.800 11.430 0.960 ;
        RECT  8.610 1.440 9.640 1.600 ;
        RECT  10.940 1.500 11.720 1.680 ;
        RECT  9.480 1.440 9.640 2.100 ;
        RECT  8.610 1.440 8.770 2.100 ;
        RECT  6.730 1.940 8.770 2.100 ;
        RECT  10.940 0.800 11.100 2.100 ;
        RECT  9.480 1.940 11.100 2.100 ;
        RECT  11.480 1.500 11.720 2.100 ;
        RECT  10.460 0.300 11.750 0.460 ;
        RECT  11.590 0.300 11.750 0.920 ;
        RECT  11.590 0.760 12.500 0.920 ;
        RECT  12.300 0.760 12.500 1.240 ;
        RECT  10.460 0.300 10.630 1.760 ;
        RECT  10.280 1.500 10.630 1.760 ;
        RECT  12.660 0.390 12.860 2.100 ;
        RECT  12.660 0.940 13.520 1.220 ;
        RECT  11.620 1.120 12.040 1.280 ;
        RECT  11.880 1.120 12.040 1.680 ;
        RECT  11.880 1.480 12.900 1.680 ;
        RECT  12.660 0.940 12.900 2.100 ;
        LAYER VTPH ;
        RECT  5.790 1.110 8.540 2.400 ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  3.310 1.090 4.120 2.400 ;
        RECT  0.000 1.200 4.120 2.400 ;
        RECT  5.790 1.140 15.600 2.400 ;
        RECT  0.000 1.210 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.090 ;
        RECT  4.120 0.000 15.600 1.110 ;
        RECT  0.000 0.000 3.310 1.140 ;
        RECT  8.540 0.000 15.600 1.140 ;
        RECT  0.500 0.000 3.310 1.200 ;
        RECT  4.120 0.000 5.790 1.210 ;
    END
END DFEQZRM8HM

MACRO DFEQZRM4HM
    CLASS CORE ;
    FOREIGN DFEQZRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.581  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 0.970 3.500 1.170 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.580 ;
        LAYER ME1 ;
        RECT  3.200 0.970 3.640 1.270 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 0.440 4.880 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.330 0.730 1.910 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.760 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.660 1.460 13.900 2.100 ;
        RECT  13.700 0.400 13.900 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  14.180 1.480 14.460 2.540 ;
        RECT  13.140 1.480 13.420 2.540 ;
        RECT  12.100 1.900 12.380 2.540 ;
        RECT  8.930 1.770 9.210 2.540 ;
        RECT  5.100 1.860 5.380 2.540 ;
        RECT  3.000 1.860 3.280 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  14.180 -0.140 14.460 0.680 ;
        RECT  13.140 -0.140 13.420 0.670 ;
        RECT  12.160 -0.140 12.320 0.600 ;
        RECT  8.930 -0.140 9.210 0.320 ;
        RECT  5.580 -0.140 6.250 0.760 ;
        RECT  3.850 -0.140 4.130 0.320 ;
        RECT  0.620 -0.140 0.900 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.330 0.380 0.600 ;
        RECT  2.190 1.060 2.660 1.220 ;
        RECT  0.100 0.330 0.260 1.940 ;
        RECT  0.900 0.760 1.060 1.540 ;
        RECT  2.190 1.060 2.440 1.540 ;
        RECT  0.100 1.380 2.440 1.540 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.060 0.330 3.360 0.490 ;
        RECT  1.060 0.330 1.470 0.540 ;
        RECT  2.070 0.650 4.340 0.810 ;
        RECT  4.060 0.650 4.340 0.990 ;
        RECT  5.040 0.380 5.200 1.380 ;
        RECT  5.040 1.180 5.930 1.380 ;
        RECT  4.340 1.220 5.930 1.380 ;
        RECT  4.340 1.220 4.620 1.730 ;
        RECT  7.010 0.300 7.570 0.610 ;
        RECT  7.370 0.300 7.570 0.660 ;
        RECT  6.620 0.420 6.810 1.420 ;
        RECT  6.620 1.140 7.780 1.420 ;
        RECT  6.090 1.260 7.780 1.420 ;
        RECT  6.090 1.260 6.250 1.780 ;
        RECT  2.600 1.540 3.920 1.700 ;
        RECT  4.780 1.540 5.700 1.700 ;
        RECT  3.560 1.540 3.920 1.740 ;
        RECT  6.410 1.580 7.810 1.740 ;
        RECT  3.760 1.540 3.920 2.100 ;
        RECT  5.540 1.540 5.700 2.100 ;
        RECT  2.600 1.540 2.760 2.080 ;
        RECT  1.620 1.800 2.760 2.080 ;
        RECT  4.780 1.540 4.940 2.100 ;
        RECT  3.760 1.940 4.940 2.100 ;
        RECT  6.410 1.580 6.570 2.100 ;
        RECT  5.540 1.940 6.570 2.100 ;
        RECT  7.850 0.360 8.130 0.640 ;
        RECT  7.970 0.360 8.130 1.280 ;
        RECT  7.970 1.120 9.660 1.280 ;
        RECT  8.010 1.060 8.290 1.780 ;
        RECT  9.700 0.620 9.980 0.960 ;
        RECT  8.670 0.800 9.980 0.960 ;
        RECT  9.820 0.620 9.980 1.760 ;
        RECT  9.800 1.480 10.000 1.760 ;
        RECT  9.370 0.300 10.300 0.460 ;
        RECT  9.370 0.300 9.540 0.640 ;
        RECT  8.290 0.480 9.540 0.640 ;
        RECT  8.290 0.480 8.450 0.900 ;
        RECT  10.140 0.300 10.300 1.100 ;
        RECT  11.150 0.620 11.430 0.960 ;
        RECT  10.940 0.800 11.430 0.960 ;
        RECT  8.610 1.440 9.640 1.600 ;
        RECT  10.940 1.500 11.720 1.680 ;
        RECT  9.480 1.440 9.640 2.100 ;
        RECT  8.610 1.440 8.770 2.100 ;
        RECT  6.730 1.940 8.770 2.100 ;
        RECT  10.940 0.800 11.100 2.100 ;
        RECT  9.480 1.940 11.100 2.100 ;
        RECT  11.480 1.500 11.720 2.100 ;
        RECT  10.460 0.300 11.750 0.460 ;
        RECT  11.590 0.300 11.750 0.920 ;
        RECT  11.590 0.760 12.500 0.920 ;
        RECT  12.300 0.760 12.500 1.240 ;
        RECT  10.460 0.300 10.630 1.760 ;
        RECT  10.280 1.500 10.630 1.760 ;
        RECT  12.660 0.390 12.860 2.100 ;
        RECT  12.660 0.940 13.520 1.220 ;
        RECT  11.620 1.120 12.040 1.280 ;
        RECT  11.880 1.120 12.040 1.680 ;
        RECT  11.880 1.480 12.900 1.680 ;
        RECT  12.660 0.940 12.900 2.100 ;
        LAYER VTPH ;
        RECT  5.790 1.110 8.540 2.400 ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  3.310 1.090 4.120 2.400 ;
        RECT  0.000 1.200 4.120 2.400 ;
        RECT  5.790 1.140 14.800 2.400 ;
        RECT  0.000 1.210 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.090 ;
        RECT  4.120 0.000 14.800 1.110 ;
        RECT  0.000 0.000 3.310 1.140 ;
        RECT  8.540 0.000 14.800 1.140 ;
        RECT  0.500 0.000 3.310 1.200 ;
        RECT  4.120 0.000 5.790 1.210 ;
    END
END DFEQZRM4HM

MACRO DFEQZRM2HM
    CLASS CORE ;
    FOREIGN DFEQZRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        ANTENNAGATEAREA 0.084  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.933  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 0.970 3.500 1.170 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.580 ;
        LAYER ME1 ;
        RECT  2.820 0.970 3.640 1.270 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 0.440 4.880 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.070  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.330 0.730 1.910 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.760 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.580 1.460 13.900 2.100 ;
        RECT  13.700 0.400 13.900 2.100 ;
        RECT  13.620 0.400 13.900 0.730 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.060 1.480 13.340 2.540 ;
        RECT  12.040 1.900 12.320 2.540 ;
        RECT  8.930 1.770 9.210 2.540 ;
        RECT  5.100 1.860 5.380 2.540 ;
        RECT  3.000 1.860 3.280 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.060 -0.140 13.340 0.670 ;
        RECT  12.100 -0.140 12.260 0.600 ;
        RECT  8.930 -0.140 9.210 0.320 ;
        RECT  5.580 -0.140 6.250 0.760 ;
        RECT  3.850 -0.140 4.130 0.320 ;
        RECT  0.620 -0.140 0.900 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.330 0.380 0.600 ;
        RECT  2.190 1.060 2.660 1.220 ;
        RECT  0.100 0.330 0.260 1.940 ;
        RECT  0.900 0.760 1.060 1.540 ;
        RECT  2.190 1.060 2.440 1.540 ;
        RECT  0.100 1.380 2.440 1.540 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.060 0.330 3.360 0.490 ;
        RECT  1.060 0.330 1.470 0.540 ;
        RECT  2.070 0.650 4.340 0.810 ;
        RECT  4.060 0.650 4.340 0.990 ;
        RECT  5.040 0.380 5.200 1.380 ;
        RECT  5.040 1.180 5.930 1.380 ;
        RECT  4.340 1.220 5.930 1.380 ;
        RECT  4.340 1.220 4.620 1.730 ;
        RECT  7.010 0.300 7.570 0.610 ;
        RECT  7.370 0.300 7.570 0.660 ;
        RECT  6.620 0.420 6.810 1.420 ;
        RECT  6.620 1.140 7.780 1.420 ;
        RECT  6.090 1.260 7.780 1.420 ;
        RECT  6.090 1.260 6.250 1.780 ;
        RECT  2.600 1.540 3.920 1.700 ;
        RECT  4.780 1.540 5.700 1.700 ;
        RECT  3.560 1.540 3.920 1.740 ;
        RECT  6.410 1.580 7.810 1.740 ;
        RECT  3.760 1.540 3.920 2.100 ;
        RECT  5.540 1.540 5.700 2.100 ;
        RECT  2.600 1.540 2.760 2.080 ;
        RECT  1.620 1.800 2.760 2.080 ;
        RECT  4.780 1.540 4.940 2.100 ;
        RECT  3.760 1.940 4.940 2.100 ;
        RECT  6.410 1.580 6.570 2.100 ;
        RECT  5.540 1.940 6.570 2.100 ;
        RECT  7.850 0.360 8.130 0.640 ;
        RECT  7.970 0.360 8.130 1.280 ;
        RECT  7.970 1.120 9.660 1.280 ;
        RECT  8.010 1.060 8.290 1.780 ;
        RECT  9.700 0.620 9.980 0.960 ;
        RECT  8.670 0.800 9.980 0.960 ;
        RECT  9.820 0.620 9.980 1.760 ;
        RECT  9.800 1.480 10.000 1.760 ;
        RECT  9.370 0.300 10.300 0.460 ;
        RECT  9.370 0.300 9.540 0.640 ;
        RECT  8.290 0.480 9.540 0.640 ;
        RECT  8.290 0.480 8.450 0.900 ;
        RECT  10.140 0.300 10.300 1.100 ;
        RECT  11.150 0.620 11.430 0.960 ;
        RECT  10.940 0.800 11.430 0.960 ;
        RECT  8.610 1.440 9.640 1.600 ;
        RECT  10.940 1.500 11.720 1.680 ;
        RECT  9.480 1.440 9.640 2.100 ;
        RECT  8.610 1.440 8.770 2.100 ;
        RECT  6.730 1.940 8.770 2.100 ;
        RECT  10.940 0.800 11.100 2.100 ;
        RECT  9.480 1.940 11.100 2.100 ;
        RECT  11.480 1.500 11.720 2.100 ;
        RECT  10.460 0.300 11.750 0.460 ;
        RECT  11.590 0.300 11.750 0.920 ;
        RECT  11.590 0.760 12.420 0.920 ;
        RECT  12.220 0.760 12.420 1.240 ;
        RECT  10.460 0.300 10.630 1.760 ;
        RECT  10.280 1.500 10.630 1.760 ;
        RECT  12.580 0.390 12.780 2.100 ;
        RECT  12.580 0.940 13.440 1.220 ;
        RECT  11.620 1.120 12.040 1.280 ;
        RECT  11.880 1.120 12.040 1.680 ;
        RECT  11.880 1.480 12.820 1.680 ;
        RECT  12.580 0.940 12.820 2.100 ;
        LAYER VTPH ;
        RECT  5.790 1.110 8.540 2.400 ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  3.310 1.090 4.120 2.400 ;
        RECT  0.000 1.200 4.120 2.400 ;
        RECT  5.790 1.140 14.000 2.400 ;
        RECT  0.000 1.210 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.090 ;
        RECT  4.120 0.000 14.000 1.110 ;
        RECT  0.000 0.000 3.310 1.140 ;
        RECT  8.540 0.000 14.000 1.140 ;
        RECT  0.500 0.000 3.310 1.200 ;
        RECT  4.120 0.000 5.790 1.210 ;
    END
END DFEQZRM2HM

MACRO DFEQZRM1HM
    CLASS CORE ;
    FOREIGN DFEQZRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        ANTENNAGATEAREA 0.071  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 8.226  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 0.970 3.500 1.170 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.580 ;
        LAYER ME1 ;
        RECT  2.820 0.970 3.640 1.270 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 0.440 4.880 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.330 0.730 1.910 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.760 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.620 1.460 13.900 1.740 ;
        RECT  13.700 0.320 13.900 1.740 ;
        RECT  13.660 0.320 13.900 0.730 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.100 1.480 13.380 2.540 ;
        RECT  12.080 1.900 12.360 2.540 ;
        RECT  8.930 1.770 9.210 2.540 ;
        RECT  5.100 1.860 5.380 2.540 ;
        RECT  3.000 1.860 3.280 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.100 -0.140 13.380 0.600 ;
        RECT  12.140 -0.140 12.300 0.600 ;
        RECT  8.930 -0.140 9.210 0.320 ;
        RECT  5.580 -0.140 6.250 0.760 ;
        RECT  3.850 -0.140 4.130 0.320 ;
        RECT  0.620 -0.140 0.900 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.330 0.380 0.600 ;
        RECT  2.190 1.060 2.610 1.220 ;
        RECT  0.100 0.330 0.260 1.940 ;
        RECT  0.900 0.760 1.060 1.540 ;
        RECT  2.190 1.060 2.350 1.540 ;
        RECT  0.100 1.380 2.350 1.540 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.060 0.330 3.360 0.490 ;
        RECT  1.060 0.330 1.470 0.540 ;
        RECT  2.070 0.650 4.340 0.810 ;
        RECT  4.060 0.650 4.340 0.990 ;
        RECT  5.040 0.380 5.200 1.380 ;
        RECT  5.040 1.180 5.930 1.380 ;
        RECT  4.340 1.220 5.930 1.380 ;
        RECT  4.340 1.220 4.620 1.730 ;
        RECT  7.010 0.300 7.570 0.610 ;
        RECT  6.620 0.420 6.810 1.420 ;
        RECT  6.620 1.140 7.780 1.420 ;
        RECT  6.090 1.260 7.780 1.420 ;
        RECT  6.090 1.260 6.250 1.780 ;
        RECT  2.600 1.540 3.920 1.700 ;
        RECT  4.780 1.540 5.700 1.700 ;
        RECT  3.560 1.540 3.920 1.740 ;
        RECT  6.410 1.580 7.810 1.740 ;
        RECT  2.600 1.540 2.760 1.910 ;
        RECT  1.580 1.750 2.760 1.910 ;
        RECT  3.760 1.540 3.920 2.100 ;
        RECT  5.540 1.540 5.700 2.100 ;
        RECT  4.780 1.540 4.940 2.100 ;
        RECT  3.760 1.940 4.940 2.100 ;
        RECT  6.410 1.580 6.570 2.100 ;
        RECT  5.540 1.940 6.570 2.100 ;
        RECT  7.850 0.300 8.130 0.610 ;
        RECT  7.970 0.300 8.130 1.280 ;
        RECT  7.970 1.120 9.660 1.280 ;
        RECT  8.010 1.060 8.290 1.780 ;
        RECT  9.700 0.620 9.980 0.960 ;
        RECT  8.670 0.800 9.980 0.960 ;
        RECT  9.820 0.620 9.980 1.760 ;
        RECT  9.800 1.480 10.000 1.760 ;
        RECT  9.370 0.300 10.300 0.460 ;
        RECT  9.370 0.300 9.540 0.640 ;
        RECT  8.290 0.480 9.540 0.640 ;
        RECT  8.290 0.480 8.450 0.900 ;
        RECT  10.140 0.300 10.300 1.100 ;
        RECT  11.150 0.620 11.430 0.960 ;
        RECT  10.940 0.800 11.430 0.960 ;
        RECT  8.610 1.440 9.640 1.600 ;
        RECT  10.940 1.500 11.720 1.680 ;
        RECT  9.480 1.440 9.640 2.100 ;
        RECT  8.610 1.440 8.770 2.100 ;
        RECT  6.730 1.940 8.770 2.100 ;
        RECT  10.940 0.800 11.100 2.100 ;
        RECT  9.480 1.940 11.100 2.100 ;
        RECT  11.480 1.500 11.720 2.100 ;
        RECT  10.460 0.300 11.750 0.460 ;
        RECT  11.590 0.300 11.750 0.920 ;
        RECT  11.590 0.760 12.460 0.920 ;
        RECT  12.260 0.760 12.460 1.240 ;
        RECT  10.460 0.300 10.630 1.760 ;
        RECT  10.280 1.500 10.630 1.760 ;
        RECT  12.620 0.320 12.820 1.740 ;
        RECT  12.620 0.940 13.480 1.220 ;
        RECT  11.620 1.120 12.040 1.280 ;
        RECT  11.880 1.120 12.040 1.680 ;
        RECT  11.880 1.480 12.860 1.680 ;
        RECT  12.620 0.940 12.860 1.740 ;
        RECT  12.580 1.480 12.860 1.740 ;
        LAYER VTPH ;
        RECT  5.790 1.110 8.540 2.400 ;
        RECT  0.000 1.140 0.500 2.400 ;
        RECT  3.310 1.090 4.120 2.400 ;
        RECT  0.000 1.200 4.120 2.400 ;
        RECT  5.790 1.140 14.000 2.400 ;
        RECT  0.000 1.210 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.090 ;
        RECT  4.120 0.000 14.000 1.110 ;
        RECT  0.000 0.000 3.310 1.140 ;
        RECT  8.540 0.000 14.000 1.140 ;
        RECT  0.500 0.000 3.310 1.200 ;
        RECT  4.120 0.000 5.790 1.210 ;
    END
END DFEQZRM1HM

MACRO DFEQRM8HM
    CLASS CORE ;
    FOREIGN DFEQRM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.270  LAYER ME1  ;
        ANTENNAGATEAREA 0.270  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 14.136  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 3.510 4.300 3.710 ;
        LAYER ME2 ;
        RECT  4.100 3.240 4.300 3.960 ;
        LAYER ME1 ;
        RECT  7.690 3.400 8.340 3.560 ;
        RECT  7.690 2.760 7.850 3.560 ;
        RECT  6.290 2.760 7.850 2.920 ;
        RECT  6.290 2.760 6.450 3.670 ;
        RECT  4.040 3.510 6.450 3.670 ;
        RECT  2.600 3.560 4.550 3.720 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 2.720 1.900 4.410 ;
        RECT  0.660 3.630 1.900 3.960 ;
        RECT  0.660 2.720 0.860 4.410 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  4.360 2.260 4.640 2.900 ;
        RECT  4.240 1.860 4.520 2.540 ;
        RECT  3.300 2.260 3.580 2.900 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  2.180 2.260 2.460 2.900 ;
        RECT  1.180 2.260 1.380 3.320 ;
        RECT  0.660 1.700 0.860 2.540 ;
        RECT  0.140 2.260 0.340 3.320 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  8.780 -0.140 9.060 0.500 ;
        RECT  4.780 -0.140 5.060 0.740 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        RECT  0.000 4.660 9.200 4.940 ;
        RECT  8.550 4.260 8.830 4.940 ;
        RECT  4.380 4.240 4.580 4.940 ;
        RECT  2.180 4.280 2.460 4.940 ;
        RECT  1.180 4.130 1.380 4.940 ;
        RECT  0.140 4.120 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.830 2.800 0.990 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.830 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 1.980 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 0.990 ;
        RECT  3.860 2.850 4.060 3.230 ;
        RECT  2.820 2.850 3.020 3.280 ;
        RECT  3.860 3.060 5.060 3.230 ;
        RECT  2.100 3.080 4.050 3.280 ;
        RECT  2.100 3.080 2.260 4.080 ;
        RECT  2.100 3.920 3.090 4.080 ;
        RECT  2.930 3.920 3.090 4.460 ;
        RECT  2.930 4.280 3.750 4.460 ;
        RECT  4.240 0.910 5.100 1.190 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  3.480 1.220 4.400 1.380 ;
        RECT  3.480 1.220 3.760 1.730 ;
        RECT  5.220 2.700 6.080 2.990 ;
        RECT  5.220 2.700 5.500 3.350 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  5.580 1.520 6.370 1.680 ;
        RECT  3.920 1.540 4.840 1.700 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.680 1.540 4.840 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.920 1.540 4.080 2.100 ;
        RECT  3.160 1.940 4.080 2.100 ;
        RECT  5.580 1.520 5.740 2.100 ;
        RECT  4.680 1.940 5.740 2.100 ;
        RECT  5.260 0.420 5.660 1.300 ;
        RECT  5.260 1.080 6.460 1.300 ;
        RECT  5.260 0.420 5.420 1.780 ;
        RECT  5.090 1.410 5.420 1.780 ;
        RECT  5.850 0.300 6.480 0.580 ;
        RECT  5.220 4.210 5.500 4.420 ;
        RECT  5.220 4.260 6.710 4.420 ;
        RECT  6.610 3.150 6.890 4.100 ;
        RECT  4.780 3.890 5.840 4.050 ;
        RECT  3.260 3.920 4.900 4.080 ;
        RECT  3.260 3.900 3.540 4.100 ;
        RECT  5.710 3.940 7.210 4.100 ;
        RECT  7.050 3.940 7.210 4.400 ;
        RECT  4.740 3.920 4.900 4.500 ;
        RECT  5.980 1.940 7.270 2.100 ;
        RECT  6.760 0.300 8.620 0.460 ;
        RECT  8.340 0.300 8.620 0.800 ;
        RECT  6.760 0.300 7.050 1.680 ;
        RECT  7.360 1.480 8.640 1.720 ;
        RECT  7.210 3.150 7.530 3.430 ;
        RECT  7.370 3.150 7.530 4.100 ;
        RECT  8.560 2.770 8.720 4.100 ;
        RECT  7.370 3.940 8.720 4.100 ;
        RECT  7.950 3.940 8.230 4.330 ;
        RECT  7.480 1.940 8.840 2.100 ;
        LAYER VTPH ;
        RECT  0.400 1.100 2.250 3.660 ;
        RECT  0.000 1.140 2.250 3.660 ;
        RECT  4.780 1.140 9.200 3.550 ;
        RECT  0.000 1.200 9.200 3.550 ;
        RECT  0.000 1.200 2.980 3.660 ;
        RECT  5.060 1.140 9.200 3.660 ;
        RECT  5.060 1.140 7.820 3.680 ;
        LAYER VTNH ;
        RECT  2.980 3.550 5.060 4.800 ;
        RECT  0.000 3.660 5.060 4.800 ;
        RECT  7.820 3.660 9.200 4.800 ;
        RECT  0.000 3.680 9.200 4.800 ;
        RECT  0.000 0.000 9.200 1.100 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  2.250 0.000 9.200 1.140 ;
        RECT  2.250 0.000 4.780 1.200 ;
    END
END DFEQRM8HM

MACRO DFEQRM4HM
    CLASS CORE ;
    FOREIGN DFEQRM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.229  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 3.450 1.100 3.650 ;
        LAYER ME2 ;
        RECT  0.900 3.240 1.100 3.960 ;
        LAYER ME1 ;
        RECT  0.800 3.450 1.310 3.750 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.150 0.780 1.600 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 3.660 2.770 3.820 ;
        RECT  2.550 3.360 2.770 3.820 ;
        RECT  0.420 3.910 2.010 4.070 ;
        RECT  1.540 3.660 2.010 4.070 ;
        RECT  0.420 3.750 0.640 4.070 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.530  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.830 3.030 7.170 3.560 ;
        RECT  6.630 4.100 6.990 4.380 ;
        RECT  6.830 3.030 6.990 4.380 ;
        RECT  6.600 3.030 7.170 3.190 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.240 3.560 6.030 3.840 ;
        RECT  4.240 3.560 4.760 3.990 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.760 1.770 8.040 2.540 ;
        RECT  3.250 2.260 3.530 2.930 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.890 -0.140 8.170 0.750 ;
        RECT  4.650 -0.140 4.930 0.540 ;
        RECT  0.610 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 8.400 4.940 ;
        RECT  7.190 4.190 7.420 4.940 ;
        RECT  6.030 4.480 6.310 4.940 ;
        RECT  3.980 4.480 4.270 4.940 ;
        RECT  0.640 4.300 0.920 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.990 ;
        RECT  0.100 0.710 1.000 0.990 ;
        RECT  0.100 0.300 0.260 2.070 ;
        RECT  0.100 1.770 0.320 2.070 ;
        RECT  1.170 0.320 1.500 0.600 ;
        RECT  1.280 0.320 1.500 1.770 ;
        RECT  1.090 1.520 1.500 1.770 ;
        RECT  0.100 2.850 0.380 3.250 ;
        RECT  0.100 3.090 2.340 3.250 ;
        RECT  2.060 3.090 2.340 3.460 ;
        RECT  0.100 2.850 0.260 4.500 ;
        RECT  0.100 4.230 0.380 4.500 ;
        RECT  1.270 2.770 3.090 2.930 ;
        RECT  2.930 2.770 3.090 4.140 ;
        RECT  2.170 3.980 3.090 4.140 ;
        RECT  2.170 3.980 2.330 4.470 ;
        RECT  1.420 4.300 2.330 4.470 ;
        RECT  1.660 0.330 1.920 0.680 ;
        RECT  1.760 0.330 1.920 2.100 ;
        RECT  3.110 1.820 3.380 2.100 ;
        RECT  1.760 1.940 3.380 2.100 ;
        RECT  3.810 3.520 3.970 4.150 ;
        RECT  3.660 3.940 3.820 4.460 ;
        RECT  2.510 4.300 3.820 4.460 ;
        RECT  3.540 1.660 4.930 1.860 ;
        RECT  2.130 0.330 4.450 0.490 ;
        RECT  4.290 0.330 4.450 0.860 ;
        RECT  5.090 0.370 5.250 0.860 ;
        RECT  4.290 0.700 5.250 0.860 ;
        RECT  2.130 0.330 2.420 1.760 ;
        RECT  2.580 0.650 4.130 0.820 ;
        RECT  3.970 0.650 4.130 1.180 ;
        RECT  3.970 1.020 5.720 1.180 ;
        RECT  5.520 1.020 5.720 1.340 ;
        RECT  2.580 0.650 2.800 1.740 ;
        RECT  5.410 0.370 6.060 0.630 ;
        RECT  3.590 1.090 3.810 1.500 ;
        RECT  3.590 1.340 5.360 1.500 ;
        RECT  5.880 0.370 6.060 1.730 ;
        RECT  5.200 1.340 5.360 1.730 ;
        RECT  5.880 1.510 6.280 1.730 ;
        RECT  5.200 1.570 6.280 1.730 ;
        RECT  4.570 3.030 6.390 3.190 ;
        RECT  6.230 3.570 6.610 3.850 ;
        RECT  6.230 3.030 6.390 4.190 ;
        RECT  5.000 4.030 6.390 4.190 ;
        RECT  6.270 0.470 6.730 0.750 ;
        RECT  6.570 0.470 6.730 2.100 ;
        RECT  6.570 1.710 6.840 2.100 ;
        RECT  5.130 1.900 6.840 2.100 ;
        RECT  6.920 0.300 7.280 0.520 ;
        RECT  6.920 0.300 7.120 1.550 ;
        RECT  7.280 0.710 7.560 1.590 ;
        RECT  7.280 1.310 8.200 1.590 ;
        RECT  7.280 0.710 7.450 1.990 ;
        RECT  7.160 1.710 7.450 1.990 ;
        RECT  4.150 2.700 8.220 2.860 ;
        RECT  7.960 2.700 8.220 3.250 ;
        RECT  4.150 2.700 4.310 3.320 ;
        RECT  3.330 3.160 4.310 3.320 ;
        RECT  3.330 3.160 3.490 3.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.760 3.660 ;
        RECT  0.000 1.200 4.590 3.660 ;
        RECT  5.820 1.210 7.040 3.660 ;
        RECT  0.000 1.260 7.040 3.660 ;
        RECT  7.940 1.140 8.400 3.660 ;
        RECT  0.000 1.270 8.400 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 8.400 4.800 ;
        RECT  0.000 0.000 8.400 1.140 ;
        RECT  2.760 0.000 7.940 1.200 ;
        RECT  4.590 0.000 7.940 1.210 ;
        RECT  4.590 0.000 5.820 1.260 ;
        RECT  7.040 0.000 7.940 1.270 ;
    END
END DFEQRM4HM

MACRO DFEQRM2HM
    CLASS CORE ;
    FOREIGN DFEQRM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.100  LAYER ME1  ;
        ANTENNAGATEAREA 0.100  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.229  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 3.450 1.100 3.650 ;
        LAYER ME2 ;
        RECT  0.900 3.240 1.100 3.960 ;
        LAYER ME1 ;
        RECT  0.800 3.450 1.310 3.750 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.150 0.780 1.600 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 3.660 2.770 3.820 ;
        RECT  2.550 3.360 2.770 3.820 ;
        RECT  0.420 3.910 2.010 4.070 ;
        RECT  1.540 3.660 2.010 4.070 ;
        RECT  0.420 3.750 0.640 4.070 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 4.040 6.450 4.380 ;
        RECT  6.240 3.030 6.450 4.380 ;
        RECT  6.120 3.030 6.450 3.350 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.167  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.240 3.560 4.760 4.010 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.260 2.260 7.540 3.270 ;
        RECT  3.250 2.260 3.530 2.930 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  4.650 -0.140 4.930 0.540 ;
        RECT  0.610 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 8.000 4.940 ;
        RECT  7.210 4.160 7.490 4.940 ;
        RECT  5.550 4.480 5.830 4.940 ;
        RECT  3.980 4.480 4.270 4.940 ;
        RECT  0.640 4.300 0.920 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.990 ;
        RECT  0.100 0.710 1.000 0.990 ;
        RECT  0.100 0.300 0.260 2.070 ;
        RECT  0.100 1.770 0.320 2.070 ;
        RECT  1.170 0.320 1.500 0.600 ;
        RECT  1.280 0.320 1.500 1.770 ;
        RECT  1.090 1.520 1.500 1.770 ;
        RECT  0.100 2.850 0.380 3.250 ;
        RECT  0.100 3.090 2.340 3.250 ;
        RECT  2.060 3.090 2.340 3.460 ;
        RECT  0.100 2.850 0.260 4.500 ;
        RECT  0.100 4.230 0.380 4.500 ;
        RECT  1.270 2.770 3.090 2.930 ;
        RECT  2.930 2.770 3.090 4.140 ;
        RECT  2.170 3.980 3.090 4.140 ;
        RECT  2.170 3.980 2.330 4.470 ;
        RECT  1.420 4.300 2.330 4.470 ;
        RECT  1.660 0.330 1.920 0.680 ;
        RECT  1.760 0.330 1.920 2.100 ;
        RECT  3.110 1.820 3.380 2.100 ;
        RECT  1.760 1.940 3.380 2.100 ;
        RECT  3.810 3.520 3.970 4.150 ;
        RECT  3.660 3.940 3.820 4.460 ;
        RECT  2.510 4.300 3.820 4.460 ;
        RECT  3.540 1.660 4.900 1.860 ;
        RECT  2.130 0.330 4.180 0.490 ;
        RECT  4.020 0.330 4.180 0.860 ;
        RECT  5.090 0.370 5.250 0.860 ;
        RECT  4.020 0.700 5.250 0.860 ;
        RECT  2.130 0.330 2.420 1.760 ;
        RECT  2.580 0.650 3.860 0.820 ;
        RECT  3.700 0.650 3.860 1.180 ;
        RECT  3.700 1.020 5.620 1.180 ;
        RECT  5.420 1.020 5.620 1.340 ;
        RECT  2.580 0.650 2.800 1.740 ;
        RECT  4.570 3.030 5.910 3.190 ;
        RECT  5.750 3.570 6.030 3.850 ;
        RECT  5.750 3.030 5.910 4.190 ;
        RECT  5.000 4.030 5.910 4.190 ;
        RECT  5.410 0.370 5.940 0.630 ;
        RECT  3.320 1.090 3.540 1.500 ;
        RECT  3.320 1.340 5.260 1.500 ;
        RECT  5.780 0.370 5.940 1.730 ;
        RECT  5.100 1.340 5.260 1.730 ;
        RECT  5.780 1.510 6.280 1.730 ;
        RECT  5.100 1.570 6.280 1.730 ;
        RECT  6.100 0.470 6.600 0.750 ;
        RECT  6.440 0.470 6.600 2.100 ;
        RECT  6.440 1.710 6.840 2.100 ;
        RECT  5.130 1.900 6.840 2.100 ;
        RECT  4.150 2.700 6.930 2.860 ;
        RECT  4.150 2.700 4.310 3.320 ;
        RECT  3.330 3.160 4.310 3.320 ;
        RECT  3.330 3.160 3.490 3.740 ;
        RECT  6.610 2.700 6.930 4.380 ;
        RECT  6.760 0.300 7.040 0.540 ;
        RECT  6.760 0.300 6.980 1.410 ;
        RECT  7.140 0.710 7.480 1.710 ;
        RECT  7.160 0.710 7.480 1.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.760 3.660 ;
        RECT  5.820 1.210 6.920 3.660 ;
        RECT  0.000 1.200 4.210 3.660 ;
        RECT  5.820 1.230 8.000 3.660 ;
        RECT  0.000 1.260 8.000 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 8.000 4.800 ;
        RECT  0.000 0.000 8.000 1.140 ;
        RECT  2.760 0.000 8.000 1.200 ;
        RECT  4.210 0.000 8.000 1.210 ;
        RECT  6.920 0.000 8.000 1.230 ;
        RECT  4.210 0.000 5.820 1.260 ;
    END
END DFEQRM2HM

MACRO DFEQRM1HM
    CLASS CORE ;
    FOREIGN DFEQRM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        ANTENNAGATEAREA 0.077  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.484  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 3.450 1.100 3.650 ;
        LAYER ME2 ;
        RECT  0.900 3.240 1.100 3.960 ;
        LAYER ME1 ;
        RECT  0.800 3.450 1.310 3.750 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.150 0.780 1.600 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 3.660 2.770 3.820 ;
        RECT  2.550 3.360 2.770 3.820 ;
        RECT  0.420 3.910 2.010 4.070 ;
        RECT  1.540 3.660 2.010 4.070 ;
        RECT  0.420 3.750 0.640 4.070 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 4.040 6.450 4.410 ;
        RECT  6.240 3.030 6.450 4.410 ;
        RECT  6.120 3.030 6.450 3.350 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.240 3.560 4.760 4.020 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.260 2.260 7.540 3.270 ;
        RECT  3.250 2.260 3.530 2.930 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  4.650 -0.140 4.930 0.540 ;
        RECT  0.610 -0.140 0.900 0.540 ;
        RECT  0.000 4.660 8.000 4.940 ;
        RECT  7.210 4.160 7.490 4.940 ;
        RECT  5.550 4.480 5.830 4.940 ;
        RECT  3.980 4.480 4.270 4.940 ;
        RECT  0.640 4.300 0.920 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.300 0.380 0.990 ;
        RECT  0.100 0.710 1.000 0.990 ;
        RECT  0.100 0.300 0.260 2.060 ;
        RECT  0.100 1.780 0.320 2.060 ;
        RECT  1.170 0.320 1.500 0.600 ;
        RECT  1.280 0.320 1.500 1.910 ;
        RECT  1.090 1.660 1.500 1.910 ;
        RECT  0.100 2.860 0.380 3.250 ;
        RECT  0.100 3.090 2.340 3.250 ;
        RECT  2.060 3.090 2.340 3.460 ;
        RECT  0.100 2.860 0.260 4.500 ;
        RECT  0.100 4.240 0.380 4.500 ;
        RECT  1.270 2.770 3.090 2.930 ;
        RECT  2.930 2.770 3.090 4.140 ;
        RECT  2.170 3.980 3.090 4.140 ;
        RECT  2.170 3.980 2.330 4.470 ;
        RECT  1.420 4.300 2.330 4.470 ;
        RECT  1.660 0.330 1.920 0.680 ;
        RECT  1.760 0.330 1.920 2.100 ;
        RECT  3.110 1.820 3.380 2.100 ;
        RECT  1.760 1.940 3.380 2.100 ;
        RECT  3.810 3.520 3.970 4.150 ;
        RECT  3.660 3.940 3.820 4.460 ;
        RECT  2.510 4.300 3.820 4.460 ;
        RECT  3.540 1.660 4.900 1.860 ;
        RECT  2.130 0.330 4.180 0.490 ;
        RECT  4.020 0.330 4.180 0.860 ;
        RECT  5.090 0.370 5.250 0.860 ;
        RECT  4.020 0.700 5.250 0.860 ;
        RECT  2.130 0.330 2.420 1.760 ;
        RECT  2.580 0.650 3.860 0.820 ;
        RECT  3.700 0.650 3.860 1.180 ;
        RECT  3.700 1.020 5.620 1.180 ;
        RECT  5.420 1.020 5.620 1.340 ;
        RECT  2.580 0.650 2.800 1.740 ;
        RECT  4.570 3.030 5.910 3.190 ;
        RECT  5.750 3.570 6.030 3.850 ;
        RECT  5.750 3.030 5.910 4.320 ;
        RECT  5.000 4.160 5.910 4.320 ;
        RECT  5.410 0.370 5.940 0.630 ;
        RECT  3.320 1.090 3.540 1.500 ;
        RECT  3.320 1.340 5.260 1.500 ;
        RECT  5.780 0.370 5.940 1.730 ;
        RECT  5.100 1.340 5.260 1.730 ;
        RECT  5.780 1.510 6.280 1.730 ;
        RECT  5.100 1.570 6.280 1.730 ;
        RECT  6.100 0.470 6.600 0.750 ;
        RECT  6.440 0.470 6.600 2.100 ;
        RECT  6.440 1.710 6.840 2.100 ;
        RECT  5.130 1.900 6.840 2.100 ;
        RECT  4.150 2.700 6.930 2.860 ;
        RECT  4.150 2.700 4.310 3.320 ;
        RECT  3.330 3.160 4.310 3.320 ;
        RECT  3.330 3.160 3.490 3.740 ;
        RECT  6.610 2.700 6.930 4.380 ;
        RECT  6.760 0.300 7.040 0.540 ;
        RECT  6.760 0.300 6.980 1.410 ;
        RECT  7.140 0.710 7.480 1.710 ;
        RECT  7.160 0.710 7.480 1.990 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.760 3.660 ;
        RECT  5.820 1.210 6.920 3.660 ;
        RECT  0.000 1.200 4.210 3.660 ;
        RECT  5.820 1.230 8.000 3.660 ;
        RECT  0.000 1.260 8.000 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 8.000 4.800 ;
        RECT  0.000 0.000 8.000 1.140 ;
        RECT  2.760 0.000 8.000 1.200 ;
        RECT  4.210 0.000 8.000 1.210 ;
        RECT  6.920 0.000 8.000 1.230 ;
        RECT  4.210 0.000 5.820 1.260 ;
    END
END DFEQRM1HM

MACRO DFEQM8HM
    CLASS CORE ;
    FOREIGN DFEQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.900 0.400 14.220 2.100 ;
        RECT  12.900 0.840 14.220 1.170 ;
        RECT  12.860 1.460 13.100 2.100 ;
        RECT  12.900 0.400 13.100 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  14.420 1.480 14.700 2.540 ;
        RECT  13.380 1.480 13.660 2.540 ;
        RECT  12.340 1.480 12.620 2.540 ;
        RECT  11.300 1.900 11.580 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  14.420 -0.140 14.700 0.680 ;
        RECT  13.380 -0.140 13.660 0.680 ;
        RECT  12.340 -0.140 12.620 0.670 ;
        RECT  11.360 -0.140 11.520 0.600 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.830 2.800 0.990 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.830 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 1.980 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 0.990 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  10.350 0.620 10.630 0.960 ;
        RECT  10.140 0.800 10.630 0.960 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.140 1.500 10.920 1.680 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  10.140 0.800 10.300 2.100 ;
        RECT  8.680 1.940 10.300 2.100 ;
        RECT  10.680 1.500 10.920 2.100 ;
        RECT  9.660 0.300 10.950 0.460 ;
        RECT  10.790 0.300 10.950 0.920 ;
        RECT  10.790 0.760 11.700 0.920 ;
        RECT  11.500 0.760 11.700 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.860 0.390 12.060 2.100 ;
        RECT  11.860 0.940 12.720 1.220 ;
        RECT  10.820 1.120 11.240 1.280 ;
        RECT  11.080 1.120 11.240 1.680 ;
        RECT  11.080 1.480 12.100 1.680 ;
        RECT  11.860 0.940 12.100 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 14.800 2.400 ;
        RECT  0.000 1.210 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 14.800 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEQM8HM

MACRO DFEQM4HM
    CLASS CORE ;
    FOREIGN DFEQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.860 1.460 13.100 2.100 ;
        RECT  12.900 0.400 13.100 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.380 1.480 13.660 2.540 ;
        RECT  12.340 1.480 12.620 2.540 ;
        RECT  11.300 1.900 11.580 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.380 -0.140 13.660 0.680 ;
        RECT  12.340 -0.140 12.620 0.670 ;
        RECT  11.360 -0.140 11.520 0.600 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.880 2.800 1.040 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.880 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 1.980 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 1.040 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  10.350 0.620 10.630 0.960 ;
        RECT  10.140 0.800 10.630 0.960 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.140 1.500 10.920 1.680 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  10.140 0.800 10.300 2.100 ;
        RECT  8.680 1.940 10.300 2.100 ;
        RECT  10.680 1.500 10.920 2.100 ;
        RECT  9.660 0.300 10.950 0.460 ;
        RECT  10.790 0.300 10.950 0.920 ;
        RECT  10.790 0.760 11.700 0.920 ;
        RECT  11.500 0.760 11.700 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.860 0.390 12.060 2.100 ;
        RECT  11.860 0.940 12.720 1.220 ;
        RECT  10.820 1.120 11.240 1.280 ;
        RECT  11.080 1.120 11.240 1.680 ;
        RECT  11.080 1.480 12.100 1.680 ;
        RECT  11.860 0.940 12.100 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 14.000 2.400 ;
        RECT  0.000 1.210 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 14.000 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEQM4HM

MACRO DFEQM2HM
    CLASS CORE ;
    FOREIGN DFEQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.820 1.460 13.100 2.100 ;
        RECT  12.900 0.400 13.100 2.100 ;
        RECT  12.820 0.400 13.100 0.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.300 1.480 12.580 2.540 ;
        RECT  11.300 1.880 11.580 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.300 -0.140 12.580 0.670 ;
        RECT  11.360 -0.140 11.520 0.600 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.880 2.800 1.040 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.880 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 1.980 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 1.040 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  10.350 0.620 10.630 0.920 ;
        RECT  10.140 0.760 10.630 0.920 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.140 1.500 10.920 1.680 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  10.140 0.760 10.300 2.100 ;
        RECT  8.680 1.940 10.300 2.100 ;
        RECT  10.680 1.500 10.920 2.100 ;
        RECT  9.660 0.300 10.950 0.460 ;
        RECT  10.790 0.300 10.950 0.920 ;
        RECT  10.790 0.760 11.660 0.920 ;
        RECT  11.460 0.760 11.660 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.820 0.390 12.020 2.100 ;
        RECT  11.820 0.940 12.680 1.220 ;
        RECT  10.820 1.120 11.240 1.280 ;
        RECT  11.080 1.120 11.240 1.680 ;
        RECT  11.080 1.480 12.060 1.680 ;
        RECT  11.820 0.940 12.060 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 13.200 2.400 ;
        RECT  0.000 1.210 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 13.200 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEQM2HM

MACRO DFEQM1HM
    CLASS CORE ;
    FOREIGN DFEQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.056  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.282  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.820 1.460 13.100 1.780 ;
        RECT  12.900 0.310 13.100 1.780 ;
        RECT  12.820 0.310 13.100 0.630 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.300 1.480 12.580 2.540 ;
        RECT  11.300 1.880 11.580 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.660 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.300 -0.140 12.580 0.580 ;
        RECT  11.360 -0.140 11.520 0.600 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.880 2.800 1.040 ;
        RECT  0.100 0.300 0.260 1.980 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.980 ;
        RECT  1.660 0.880 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.710 0.300 2.460 0.670 ;
        RECT  1.710 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 1.040 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.340 3.320 1.500 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.340 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.340 2.140 1.940 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  10.350 0.620 10.630 0.920 ;
        RECT  10.140 0.760 10.630 0.920 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.140 1.500 10.920 1.680 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  10.140 0.760 10.300 2.100 ;
        RECT  8.680 1.940 10.300 2.100 ;
        RECT  10.680 1.500 10.920 2.100 ;
        RECT  9.660 0.300 10.950 0.460 ;
        RECT  10.790 0.300 10.950 0.920 ;
        RECT  10.790 0.760 11.660 0.920 ;
        RECT  11.460 0.760 11.660 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.820 0.300 12.020 1.780 ;
        RECT  11.820 0.940 12.680 1.220 ;
        RECT  10.820 1.120 11.240 1.280 ;
        RECT  11.080 1.120 11.240 1.680 ;
        RECT  11.080 1.480 12.060 1.680 ;
        RECT  11.820 0.940 12.060 1.780 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 13.200 2.400 ;
        RECT  0.000 1.210 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 13.200 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEQM1HM

MACRO DFEM8HM
    CLASS CORE ;
    FOREIGN DFEM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.166  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.060 1.380 15.620 1.600 ;
        RECT  15.300 0.400 15.620 1.600 ;
        RECT  14.140 1.300 15.620 1.600 ;
        RECT  14.140 0.400 14.340 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.540 0.370 17.740 2.100 ;
        RECT  16.500 0.900 17.740 1.160 ;
        RECT  16.500 0.370 16.700 2.100 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.400 2.540 ;
        RECT  18.060 1.480 18.260 2.540 ;
        RECT  17.020 1.480 17.220 2.540 ;
        RECT  15.900 2.080 16.180 2.540 ;
        RECT  14.700 2.080 14.980 2.540 ;
        RECT  13.500 2.080 13.780 2.540 ;
        RECT  12.300 2.080 12.580 2.540 ;
        RECT  11.240 1.840 11.440 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.400 0.140 ;
        RECT  18.060 -0.140 18.260 0.650 ;
        RECT  17.020 -0.140 17.220 0.650 ;
        RECT  15.900 -0.140 16.180 0.680 ;
        RECT  14.700 -0.140 14.980 0.680 ;
        RECT  13.500 -0.140 13.780 0.670 ;
        RECT  12.480 -0.140 12.640 0.600 ;
        RECT  10.960 -0.140 11.240 0.320 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.830 2.800 0.990 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.830 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 1.980 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 0.990 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  9.660 0.300 10.800 0.460 ;
        RECT  11.400 0.300 12.320 0.460 ;
        RECT  10.640 0.300 10.800 0.640 ;
        RECT  11.400 0.300 11.560 0.640 ;
        RECT  10.640 0.480 11.560 0.640 ;
        RECT  12.160 0.300 12.320 0.920 ;
        RECT  12.160 0.760 12.620 0.920 ;
        RECT  12.420 0.760 12.620 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  12.980 0.940 13.880 1.220 ;
        RECT  10.950 1.120 12.260 1.290 ;
        RECT  12.100 1.120 12.260 1.600 ;
        RECT  12.980 0.390 13.180 1.600 ;
        RECT  12.100 1.400 13.180 1.600 ;
        RECT  10.200 0.620 10.480 1.720 ;
        RECT  11.720 0.620 12.000 0.960 ;
        RECT  10.200 0.800 12.000 0.960 ;
        RECT  10.200 0.800 10.510 1.720 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.140 1.480 11.940 1.660 ;
        RECT  10.140 1.480 10.960 1.720 ;
        RECT  11.780 1.480 11.940 1.920 ;
        RECT  16.040 0.880 16.240 1.920 ;
        RECT  11.780 1.760 16.240 1.920 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  10.140 1.360 10.440 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  8.680 1.940 10.440 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  12.690 1.080 15.910 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 18.400 2.400 ;
        RECT  0.000 1.210 18.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.400 1.080 ;
        RECT  0.000 0.000 12.690 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 12.690 1.140 ;
        RECT  15.910 0.000 18.400 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEM8HM

MACRO DFEM4HM
    CLASS CORE ;
    FOREIGN DFEM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.583  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.020 1.380 13.540 1.600 ;
        RECT  13.100 0.840 13.540 1.600 ;
        RECT  13.100 0.400 13.500 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.260 0.810 14.800 1.160 ;
        RECT  14.260 0.370 14.460 2.100 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.780 1.480 14.980 2.540 ;
        RECT  13.660 2.080 13.940 2.540 ;
        RECT  12.460 2.080 12.740 2.540 ;
        RECT  11.260 2.080 11.540 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.780 -0.140 14.980 0.650 ;
        RECT  13.660 -0.140 13.940 0.680 ;
        RECT  12.460 -0.140 12.740 0.670 ;
        RECT  10.960 -0.140 11.240 0.320 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.830 2.800 0.990 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.830 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 1.980 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 0.990 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  9.660 0.300 10.800 0.460 ;
        RECT  10.640 0.300 10.800 0.920 ;
        RECT  10.640 0.760 11.700 0.920 ;
        RECT  11.500 0.760 11.700 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.940 0.940 12.840 1.220 ;
        RECT  10.890 1.120 11.250 1.290 ;
        RECT  11.060 1.120 11.250 1.600 ;
        RECT  11.940 0.390 12.140 1.600 ;
        RECT  11.060 1.400 12.140 1.600 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.200 0.620 10.480 1.920 ;
        RECT  13.800 0.880 14.000 1.920 ;
        RECT  10.140 1.760 14.000 1.920 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  10.140 1.360 10.390 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  8.680 1.940 10.390 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  11.650 1.080 13.670 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 15.200 2.400 ;
        RECT  0.000 1.210 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 1.080 ;
        RECT  0.000 0.000 11.650 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 11.650 1.140 ;
        RECT  13.670 0.000 15.200 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEM4HM

MACRO DFEM2HM
    CLASS CORE ;
    FOREIGN DFEM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.730 1.100 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.730 0.700 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.445  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.340 1.380 12.700 1.600 ;
        RECT  12.380 0.400 12.700 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.401  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.540 0.840 13.900 1.160 ;
        RECT  13.540 0.370 13.740 2.100 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  12.940 2.080 13.220 2.540 ;
        RECT  11.260 2.080 11.540 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.770 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  12.940 -0.140 13.220 0.680 ;
        RECT  10.960 -0.140 11.240 0.500 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.660 -0.140 0.860 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.320 1.500 0.520 ;
        RECT  1.340 0.320 1.500 1.730 ;
        RECT  0.100 0.300 0.380 0.570 ;
        RECT  1.660 0.830 2.800 0.990 ;
        RECT  0.100 0.300 0.260 1.940 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.940 ;
        RECT  1.660 0.830 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.700 0.300 2.410 0.670 ;
        RECT  1.700 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 0.990 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.450 3.320 1.610 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.450 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.450 2.140 2.050 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  9.660 0.300 10.800 0.460 ;
        RECT  10.640 0.300 10.800 0.920 ;
        RECT  10.640 0.760 11.700 0.920 ;
        RECT  11.500 0.760 11.700 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.860 0.390 12.100 1.600 ;
        RECT  11.860 0.940 12.180 1.220 ;
        RECT  10.890 1.120 11.250 1.290 ;
        RECT  11.060 1.120 11.250 1.600 ;
        RECT  11.860 0.940 12.140 1.600 ;
        RECT  11.060 1.400 12.140 1.600 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.200 0.620 10.480 1.920 ;
        RECT  13.080 0.880 13.280 1.920 ;
        RECT  10.140 1.760 13.280 1.920 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  10.140 1.440 10.390 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  8.680 1.940 10.390 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  11.650 1.080 12.950 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 14.000 2.400 ;
        RECT  0.000 1.210 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 11.650 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 11.650 1.140 ;
        RECT  12.950 0.000 14.000 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEM2HM

MACRO DFEM1HM
    CLASS CORE ;
    FOREIGN DFEM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.440 4.080 1.060 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.730 1.180 1.220 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.750 0.740 1.220 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.318  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.340 1.380 12.700 1.600 ;
        RECT  12.380 0.310 12.700 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.282  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.540 0.840 13.900 1.160 ;
        RECT  13.540 0.310 13.740 1.840 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  12.940 2.080 13.220 2.540 ;
        RECT  11.260 2.080 11.540 2.540 ;
        RECT  8.130 1.770 8.410 2.540 ;
        RECT  4.300 1.860 4.580 2.540 ;
        RECT  2.800 1.590 3.000 2.540 ;
        RECT  0.660 1.700 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  12.940 -0.140 13.220 0.590 ;
        RECT  11.230 -0.140 11.510 0.500 ;
        RECT  8.130 -0.140 8.410 0.320 ;
        RECT  4.780 -0.140 5.450 0.760 ;
        RECT  3.100 -0.140 3.380 0.320 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.140 0.340 1.500 0.540 ;
        RECT  1.340 0.340 1.500 1.730 ;
        RECT  0.100 0.300 0.370 0.590 ;
        RECT  1.660 0.830 2.800 0.990 ;
        RECT  0.100 0.300 0.260 1.980 ;
        RECT  0.100 1.380 1.180 1.540 ;
        RECT  1.020 1.380 1.180 2.100 ;
        RECT  0.100 1.380 0.340 1.980 ;
        RECT  1.660 0.830 1.820 2.100 ;
        RECT  1.020 1.940 1.820 2.100 ;
        RECT  1.740 0.300 2.410 0.670 ;
        RECT  1.740 0.510 3.480 0.670 ;
        RECT  3.200 0.510 3.480 0.990 ;
        RECT  4.240 0.380 4.400 1.380 ;
        RECT  4.240 1.180 5.130 1.380 ;
        RECT  3.540 1.220 5.130 1.380 ;
        RECT  3.540 1.220 3.820 1.730 ;
        RECT  6.210 0.300 6.770 0.610 ;
        RECT  6.570 0.300 6.770 0.660 ;
        RECT  5.820 0.420 6.010 1.420 ;
        RECT  5.820 1.140 6.980 1.420 ;
        RECT  5.290 1.260 6.980 1.420 ;
        RECT  5.290 1.260 5.450 1.780 ;
        RECT  1.980 1.270 3.320 1.430 ;
        RECT  3.980 1.540 4.900 1.700 ;
        RECT  5.610 1.580 7.010 1.740 ;
        RECT  3.160 1.270 3.320 2.100 ;
        RECT  4.740 1.540 4.900 2.100 ;
        RECT  1.980 1.270 2.140 1.940 ;
        RECT  3.980 1.540 4.140 2.100 ;
        RECT  3.160 1.940 4.140 2.100 ;
        RECT  5.610 1.580 5.770 2.100 ;
        RECT  4.740 1.940 5.770 2.100 ;
        RECT  7.050 0.360 7.330 0.640 ;
        RECT  7.170 0.360 7.330 1.280 ;
        RECT  7.170 1.120 8.860 1.280 ;
        RECT  7.210 1.060 7.490 1.780 ;
        RECT  8.900 0.620 9.180 0.960 ;
        RECT  7.870 0.800 9.180 0.960 ;
        RECT  9.020 0.620 9.180 1.760 ;
        RECT  9.000 1.480 9.200 1.760 ;
        RECT  8.570 0.300 9.500 0.460 ;
        RECT  8.570 0.300 8.740 0.640 ;
        RECT  7.490 0.480 8.740 0.640 ;
        RECT  7.490 0.480 7.650 0.900 ;
        RECT  9.340 0.300 9.500 1.100 ;
        RECT  9.660 0.300 10.800 0.460 ;
        RECT  10.640 0.300 10.800 0.920 ;
        RECT  10.640 0.760 11.700 0.920 ;
        RECT  11.500 0.760 11.700 1.240 ;
        RECT  9.660 0.300 9.830 1.760 ;
        RECT  9.480 1.500 9.830 1.760 ;
        RECT  11.860 0.350 12.100 1.600 ;
        RECT  11.860 0.940 12.180 1.220 ;
        RECT  10.890 1.120 11.250 1.290 ;
        RECT  11.060 1.120 11.250 1.600 ;
        RECT  11.860 0.940 12.140 1.600 ;
        RECT  11.060 1.400 12.140 1.600 ;
        RECT  10.200 0.620 10.480 1.920 ;
        RECT  7.810 1.440 8.840 1.600 ;
        RECT  10.140 1.550 10.900 1.920 ;
        RECT  13.080 0.880 13.280 1.920 ;
        RECT  10.140 1.760 13.280 1.920 ;
        RECT  8.680 1.440 8.840 2.100 ;
        RECT  10.140 1.440 10.390 2.100 ;
        RECT  7.810 1.440 7.970 2.100 ;
        RECT  5.930 1.940 7.970 2.100 ;
        RECT  8.680 1.940 10.390 2.100 ;
        LAYER VTPH ;
        RECT  4.990 1.110 7.740 2.400 ;
        RECT  11.650 1.080 12.950 2.400 ;
        RECT  0.500 1.110 2.340 2.400 ;
        RECT  0.000 1.140 2.340 2.400 ;
        RECT  4.990 1.140 14.000 2.400 ;
        RECT  0.000 1.210 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.080 ;
        RECT  0.000 0.000 11.650 1.110 ;
        RECT  0.000 0.000 0.500 1.140 ;
        RECT  7.740 0.000 11.650 1.140 ;
        RECT  12.950 0.000 14.000 1.140 ;
        RECT  2.340 0.000 4.990 1.210 ;
    END
END DFEM1HM

MACRO DFCRSM8HM
    CLASS CORE ;
    FOREIGN DFCRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.178  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.128  LAYER ME1  ;
        ANTENNAGATEAREA 0.128  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.564  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.514  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.074  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.510 1.440 15.250 1.600 ;
        RECT  15.050 0.400 15.250 1.600 ;
        RECT  14.010 0.400 14.300 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.927  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  17.130 0.370 17.330 2.080 ;
        RECT  16.090 0.840 17.330 1.200 ;
        RECT  16.090 0.370 16.290 2.080 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.312  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.370 0.770 12.250 0.930 ;
        RECT  11.370 0.300 11.530 0.930 ;
        RECT  9.880 0.300 11.530 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 18.000 2.540 ;
        RECT  17.650 1.430 17.850 2.540 ;
        RECT  16.610 1.430 16.810 2.540 ;
        RECT  15.420 2.080 15.700 2.540 ;
        RECT  14.210 2.080 14.490 2.540 ;
        RECT  13.010 2.080 13.290 2.540 ;
        RECT  11.690 2.080 11.970 2.540 ;
        RECT  10.430 2.080 10.710 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 18.000 0.140 ;
        RECT  17.650 -0.140 17.850 0.650 ;
        RECT  16.610 -0.140 16.810 0.650 ;
        RECT  15.570 -0.140 15.770 0.680 ;
        RECT  14.530 -0.140 14.730 0.680 ;
        RECT  13.450 -0.140 13.730 0.500 ;
        RECT  12.170 -0.140 12.370 0.560 ;
        RECT  11.690 -0.140 11.890 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.420 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.140 0.390 0.340 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.140 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 1.860 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  11.050 0.850 11.210 1.280 ;
        RECT  12.830 1.000 13.030 1.280 ;
        RECT  11.050 1.120 13.030 1.280 ;
        RECT  13.030 0.300 13.190 0.820 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.890 1.140 ;
        RECT  13.190 0.660 13.490 1.200 ;
        RECT  10.730 0.980 10.890 1.600 ;
        RECT  13.190 0.660 13.350 1.600 ;
        RECT  10.730 1.440 13.350 1.600 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 10.570 1.660 ;
        RECT  10.410 1.500 10.570 1.920 ;
        RECT  15.710 0.970 15.910 1.920 ;
        RECT  10.410 1.760 15.910 1.920 ;
        LAYER VTPH ;
        RECT  10.750 1.080 15.590 2.400 ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 18.000 2.400 ;
        RECT  0.000 1.150 18.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 18.000 1.080 ;
        RECT  0.000 0.000 10.750 1.140 ;
        RECT  15.590 0.000 18.000 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCRSM8HM

MACRO DFCRSM4HM
    CLASS CORE ;
    FOREIGN DFCRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.514  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        ANTENNAGATEAREA 0.131  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.498  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.778  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.543  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.510 1.440 14.300 1.600 ;
        RECT  14.010 0.400 14.300 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.050 0.840 15.560 1.200 ;
        RECT  15.050 0.370 15.250 2.080 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.317  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.370 0.770 12.250 0.930 ;
        RECT  11.370 0.300 11.530 0.930 ;
        RECT  9.880 0.300 11.530 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.000 2.540 ;
        RECT  15.570 1.430 15.770 2.540 ;
        RECT  14.210 2.080 14.490 2.540 ;
        RECT  13.010 2.080 13.290 2.540 ;
        RECT  11.690 2.080 11.970 2.540 ;
        RECT  10.430 2.080 10.710 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.000 0.140 ;
        RECT  15.570 -0.140 15.770 0.650 ;
        RECT  14.530 -0.140 14.730 0.680 ;
        RECT  13.450 -0.140 13.730 0.500 ;
        RECT  12.170 -0.140 12.370 0.560 ;
        RECT  11.690 -0.140 11.890 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.420 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.140 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 2.020 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  11.050 0.850 11.210 1.280 ;
        RECT  12.830 1.000 13.030 1.280 ;
        RECT  11.050 1.120 13.030 1.280 ;
        RECT  13.030 0.300 13.190 0.820 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.890 1.140 ;
        RECT  13.190 0.660 13.490 1.200 ;
        RECT  10.730 0.980 10.890 1.600 ;
        RECT  13.190 0.660 13.350 1.600 ;
        RECT  10.730 1.440 13.350 1.600 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 10.570 1.660 ;
        RECT  10.410 1.500 10.570 1.920 ;
        RECT  14.670 0.970 14.870 1.920 ;
        RECT  10.410 1.760 14.870 1.920 ;
        LAYER VTPH ;
        RECT  10.750 1.080 14.190 2.400 ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 16.000 2.400 ;
        RECT  0.000 1.150 16.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.000 1.080 ;
        RECT  0.000 0.000 10.750 1.140 ;
        RECT  14.190 0.000 16.000 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCRSM4HM

MACRO DFCRSM2HM
    CLASS CORE ;
    FOREIGN DFCRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.778  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.345  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER ME1  ;
        ANTENNAGATEAREA 0.198  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.469  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.362  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.030 1.300 12.360 1.600 ;
        RECT  12.110 0.400 12.310 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.240 0.370 13.500 2.080 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.178  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.050 0.920 11.530 1.200 ;
        RECT  11.050 0.300 11.210 1.200 ;
        RECT  9.880 0.300 11.210 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.640 2.080 12.920 2.540 ;
        RECT  11.630 2.080 11.910 2.540 ;
        RECT  10.430 2.080 10.710 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.720 -0.140 12.920 0.680 ;
        RECT  11.440 -0.140 11.640 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.420 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.140 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 2.020 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.890 1.140 ;
        RECT  11.690 0.880 11.950 1.160 ;
        RECT  10.730 0.980 10.890 1.600 ;
        RECT  11.690 0.880 11.850 1.600 ;
        RECT  10.730 1.440 11.850 1.600 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 10.570 1.660 ;
        RECT  10.410 1.500 10.570 1.920 ;
        RECT  12.860 0.970 13.060 1.920 ;
        RECT  10.410 1.760 13.060 1.920 ;
        LAYER VTPH ;
        RECT  10.750 1.080 12.540 2.400 ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 13.600 2.400 ;
        RECT  0.000 1.150 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.080 ;
        RECT  0.000 0.000 10.750 1.140 ;
        RECT  12.540 0.000 13.600 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCRSM2HM

MACRO DFCRSM1HM
    CLASS CORE ;
    FOREIGN DFCRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        ANTENNAGATEAREA 0.067  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.810  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        ANTENNAGATEAREA 0.094  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.285  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.030 1.300 12.360 1.600 ;
        RECT  12.110 0.370 12.310 1.600 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.240 0.370 13.500 1.800 ;
        END
    END QB
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.103  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.050 0.920 11.530 1.200 ;
        RECT  11.050 0.300 11.210 1.200 ;
        RECT  9.880 0.300 11.210 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  12.640 2.080 12.920 2.540 ;
        RECT  11.630 2.080 11.910 2.540 ;
        RECT  10.430 2.080 10.710 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.720 -0.140 12.920 0.650 ;
        RECT  11.440 -0.140 11.640 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.550 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.100 0.300 0.380 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.100 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 2.080 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.890 1.140 ;
        RECT  11.690 0.880 11.950 1.160 ;
        RECT  10.730 0.980 10.890 1.600 ;
        RECT  11.690 0.880 11.850 1.600 ;
        RECT  10.730 1.440 11.850 1.600 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 10.570 1.660 ;
        RECT  10.410 1.500 10.570 1.920 ;
        RECT  12.860 0.970 13.060 1.920 ;
        RECT  10.410 1.760 13.060 1.920 ;
        LAYER VTPH ;
        RECT  10.750 1.080 12.540 2.400 ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 13.600 2.400 ;
        RECT  0.000 1.150 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.080 ;
        RECT  0.000 0.000 10.750 1.140 ;
        RECT  12.540 0.000 13.600 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCRSM1HM

MACRO DFCQRSM8HM
    CLASS CORE ;
    FOREIGN DFCQRSM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.178  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.128  LAYER ME1  ;
        ANTENNAGATEAREA 0.128  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.564  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.041  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.510 1.500 15.250 1.660 ;
        RECT  15.050 0.400 15.250 1.660 ;
        RECT  14.790 1.500 15.110 2.100 ;
        RECT  14.010 0.400 14.300 1.660 ;
        RECT  13.580 1.500 13.900 2.100 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.312  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.370 0.770 12.250 0.930 ;
        RECT  11.370 0.300 11.530 0.930 ;
        RECT  9.880 0.300 11.530 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.514  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 16.000 2.540 ;
        RECT  15.420 1.440 15.700 2.540 ;
        RECT  14.210 1.900 14.490 2.540 ;
        RECT  13.010 1.900 13.290 2.540 ;
        RECT  11.690 1.900 11.970 2.540 ;
        RECT  10.430 2.080 10.710 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 16.000 0.140 ;
        RECT  15.570 -0.140 15.770 0.680 ;
        RECT  14.530 -0.140 14.730 0.680 ;
        RECT  13.450 -0.140 13.730 0.500 ;
        RECT  12.170 -0.140 12.370 0.560 ;
        RECT  11.690 -0.140 11.890 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.420 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.140 0.390 0.340 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.140 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 1.860 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 9.830 1.660 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  11.050 0.850 11.210 1.280 ;
        RECT  12.830 1.000 13.030 1.280 ;
        RECT  11.050 1.120 13.030 1.280 ;
        RECT  13.030 0.300 13.190 0.820 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.890 1.140 ;
        RECT  13.190 0.660 13.490 1.200 ;
        RECT  10.730 0.980 10.890 1.680 ;
        RECT  13.190 0.660 13.350 1.680 ;
        RECT  10.730 1.520 13.350 1.680 ;
        RECT  11.040 1.520 11.360 2.100 ;
        RECT  12.270 1.520 12.590 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 16.000 2.400 ;
        RECT  0.000 1.150 16.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 16.000 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCQRSM8HM

MACRO DFCQRSM4HM
    CLASS CORE ;
    FOREIGN DFCQRSM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.131  LAYER ME1  ;
        ANTENNAGATEAREA 0.131  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.498  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.778  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.170 1.520 13.960 1.680 ;
        RECT  13.670 0.400 13.960 1.680 ;
        RECT  13.260 1.520 13.560 2.100 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.317  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.000 0.770 11.910 0.930 ;
        RECT  11.000 0.300 11.160 0.930 ;
        RECT  9.880 0.300 11.160 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.514  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.800 2.540 ;
        RECT  13.870 1.900 14.150 2.540 ;
        RECT  12.670 1.890 12.950 2.540 ;
        RECT  11.550 1.890 11.830 2.540 ;
        RECT  10.430 2.080 10.710 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.800 0.140 ;
        RECT  14.190 -0.140 14.390 0.680 ;
        RECT  13.110 -0.140 13.390 0.500 ;
        RECT  11.830 -0.140 12.030 0.560 ;
        RECT  11.350 -0.140 11.550 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.420 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.140 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 2.020 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 9.830 1.660 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  10.680 0.850 10.840 1.280 ;
        RECT  12.490 1.000 12.690 1.280 ;
        RECT  10.680 1.120 12.690 1.280 ;
        RECT  12.690 0.300 12.850 0.820 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.520 1.140 ;
        RECT  12.850 0.660 13.150 1.200 ;
        RECT  10.360 0.980 10.520 1.700 ;
        RECT  12.850 0.660 13.010 1.700 ;
        RECT  10.360 1.540 13.010 1.700 ;
        RECT  10.980 1.540 11.280 2.100 ;
        RECT  12.100 1.540 12.400 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 14.800 2.400 ;
        RECT  0.000 1.150 14.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.800 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCQRSM4HM

MACRO DFCQRSM2HM
    CLASS CORE ;
    FOREIGN DFCQRSM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        ANTENNAGATEAREA 0.079  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.778  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.137  LAYER ME1  ;
        ANTENNAGATEAREA 0.137  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.345  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.373  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.030 1.300 12.360 1.690 ;
        RECT  12.110 0.400 12.310 1.690 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.178  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.170 0.920 11.530 1.200 ;
        RECT  11.170 0.300 11.330 1.200 ;
        RECT  9.880 0.300 11.330 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER ME1  ;
        ANTENNAGATEAREA 0.198  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.469  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.640 1.510 12.920 2.540 ;
        RECT  11.630 2.080 11.910 2.540 ;
        RECT  10.430 1.430 10.690 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.630 -0.140 12.830 0.680 ;
        RECT  11.490 -0.140 11.690 0.560 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.420 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.140 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 2.020 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.830 1.660 ;
        RECT  8.250 1.500 9.830 1.660 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 11.010 1.140 ;
        RECT  11.690 0.880 11.950 1.160 ;
        RECT  10.850 0.980 11.010 1.680 ;
        RECT  11.690 0.880 11.850 1.680 ;
        RECT  10.850 1.520 11.850 1.680 ;
        RECT  11.000 1.520 11.340 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 13.200 2.400 ;
        RECT  0.000 1.150 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCQRSM2HM

MACRO DFCQRSM1HM
    CLASS CORE ;
    FOREIGN DFCQRSM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        ANTENNAGATEAREA 0.067  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.810  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.080 0.300 1.280 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.990 0.590 1.380 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        ANTENNAGATEAREA 0.094  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.100 2.700 1.300 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.360 1.080 2.960 1.360 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.309  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.030 1.300 12.360 1.770 ;
        RECT  12.110 0.370 12.310 1.770 ;
        END
    END Q
    PIN RB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.103  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.130 0.920 11.530 1.200 ;
        RECT  11.130 0.300 11.290 1.200 ;
        RECT  9.880 0.300 11.290 0.460 ;
        RECT  9.120 0.660 10.040 0.820 ;
        RECT  9.880 0.300 10.040 0.820 ;
        RECT  9.120 0.300 9.280 0.820 ;
        RECT  6.360 0.300 9.280 0.460 ;
        RECT  4.860 1.120 6.520 1.280 ;
        RECT  6.360 0.300 6.520 1.280 ;
        RECT  4.860 1.060 5.560 1.280 ;
        RECT  5.240 0.840 5.560 1.280 ;
        RECT  4.860 1.060 5.150 1.370 ;
        END
    END RB
    PIN SB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        ANTENNAGATEAREA 0.144  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.670 0.940 8.870 1.140 ;
        LAYER ME2 ;
        RECT  8.500 0.840 8.870 1.560 ;
        LAYER ME1 ;
        RECT  8.570 0.980 9.170 1.280 ;
        RECT  8.570 0.940 9.000 1.280 ;
        END
    END SB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.640 1.560 12.920 2.540 ;
        RECT  11.630 2.080 11.910 2.540 ;
        RECT  10.430 1.510 10.650 2.540 ;
        RECT  6.220 2.080 6.500 2.540 ;
        RECT  1.660 1.690 1.860 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.630 -0.140 12.830 0.650 ;
        RECT  11.450 -0.140 11.640 0.610 ;
        RECT  9.440 -0.140 9.720 0.500 ;
        RECT  3.830 -0.140 4.110 0.320 ;
        RECT  2.140 -0.140 2.300 0.600 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.530 1.480 4.290 1.760 ;
        RECT  2.880 0.620 3.280 0.780 ;
        RECT  4.590 0.620 4.980 0.890 ;
        RECT  3.120 0.800 4.730 0.960 ;
        RECT  3.120 0.620 3.280 1.710 ;
        RECT  2.550 1.530 3.280 1.710 ;
        RECT  1.060 0.300 1.980 0.460 ;
        RECT  2.460 0.300 3.660 0.460 ;
        RECT  4.270 0.300 6.200 0.460 ;
        RECT  3.500 0.300 3.660 0.640 ;
        RECT  4.270 0.300 4.430 0.640 ;
        RECT  3.500 0.480 4.430 0.640 ;
        RECT  0.100 0.300 0.380 0.830 ;
        RECT  1.820 0.300 1.980 0.920 ;
        RECT  1.060 0.300 1.220 0.830 ;
        RECT  0.100 0.660 1.220 0.830 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.820 0.760 2.620 0.920 ;
        RECT  5.920 0.300 6.200 0.920 ;
        RECT  0.800 0.660 1.000 1.700 ;
        RECT  0.100 1.540 1.000 1.700 ;
        RECT  0.100 1.540 0.380 2.080 ;
        RECT  1.380 0.620 1.660 0.840 ;
        RECT  1.380 0.620 1.540 1.520 ;
        RECT  1.180 1.340 2.180 1.520 ;
        RECT  5.900 1.760 7.240 1.920 ;
        RECT  2.020 1.340 2.180 2.100 ;
        RECT  1.180 1.340 1.380 2.080 ;
        RECT  5.900 1.760 6.060 2.100 ;
        RECT  2.020 1.940 6.060 2.100 ;
        RECT  3.680 1.120 4.650 1.280 ;
        RECT  6.700 0.620 6.980 1.600 ;
        RECT  6.700 1.390 7.630 1.600 ;
        RECT  5.460 1.440 7.630 1.600 ;
        RECT  4.490 1.120 4.650 1.780 ;
        RECT  7.410 1.390 7.630 1.770 ;
        RECT  5.460 1.440 5.740 1.780 ;
        RECT  4.490 1.620 5.740 1.780 ;
        RECT  7.870 0.620 8.890 0.780 ;
        RECT  7.870 0.620 8.410 0.870 ;
        RECT  8.250 0.620 8.410 1.660 ;
        RECT  8.250 1.440 8.750 1.660 ;
        RECT  9.550 1.450 9.870 1.660 ;
        RECT  8.250 1.500 9.870 1.660 ;
        RECT  7.310 0.620 7.590 1.190 ;
        RECT  7.310 1.030 8.090 1.190 ;
        RECT  7.930 1.030 8.090 1.980 ;
        RECT  7.930 1.820 10.250 1.980 ;
        RECT  9.830 1.820 10.250 2.000 ;
        RECT  10.200 0.620 10.480 1.140 ;
        RECT  9.360 0.980 10.970 1.140 ;
        RECT  11.690 0.880 11.950 1.160 ;
        RECT  10.810 0.980 10.970 1.700 ;
        RECT  11.690 0.880 11.850 1.700 ;
        RECT  10.810 1.540 11.850 1.700 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.340 2.400 ;
        RECT  8.320 1.140 13.200 2.400 ;
        RECT  0.000 1.150 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.140 ;
        RECT  6.340 0.000 8.320 1.150 ;
    END
END DFCQRSM1HM

MACRO DFCQM8HM
    CLASS CORE ;
    FOREIGN DFCQM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        ANTENNAGATEAREA 0.118  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.793  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.280 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.610 0.850 10.880 2.100 ;
        RECT  10.670 0.380 10.880 2.100 ;
        RECT  9.610 0.850 10.880 1.100 ;
        RECT  9.610 0.390 9.810 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.190 1.440 11.350 2.540 ;
        RECT  10.150 1.410 10.310 2.540 ;
        RECT  9.040 1.450 9.240 2.540 ;
        RECT  7.950 1.460 8.150 2.540 ;
        RECT  6.830 1.520 7.110 2.540 ;
        RECT  3.780 2.000 3.980 2.540 ;
        RECT  1.780 1.790 1.980 2.540 ;
        RECT  0.660 2.060 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.170 -0.140 11.370 0.660 ;
        RECT  10.130 -0.140 10.340 0.610 ;
        RECT  9.090 -0.140 9.290 0.610 ;
        RECT  8.110 -0.140 8.270 0.630 ;
        RECT  6.590 -0.140 6.870 0.320 ;
        RECT  3.860 -0.140 4.140 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.120 1.120 4.400 1.340 ;
        RECT  3.060 1.290 4.280 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.620 0.620 4.910 0.950 ;
        RECT  3.640 0.800 4.720 0.960 ;
        RECT  3.640 0.800 3.920 1.100 ;
        RECT  4.560 0.800 4.720 1.780 ;
        RECT  4.500 1.500 4.780 1.780 ;
        RECT  1.340 0.620 1.620 1.610 ;
        RECT  1.340 1.440 2.300 1.610 ;
        RECT  1.260 1.500 1.500 1.820 ;
        RECT  3.440 1.680 4.340 1.840 ;
        RECT  2.140 1.440 2.300 2.090 ;
        RECT  4.180 1.680 4.340 2.100 ;
        RECT  3.440 1.680 3.600 2.090 ;
        RECT  2.140 1.930 3.600 2.090 ;
        RECT  4.180 1.940 5.190 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.580 0.460 ;
        RECT  4.300 0.300 5.910 0.460 ;
        RECT  3.400 0.300 3.580 0.640 ;
        RECT  4.300 0.300 4.460 0.640 ;
        RECT  3.400 0.480 4.460 0.640 ;
        RECT  0.140 0.450 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.750 0.300 5.910 1.700 ;
        RECT  0.800 0.750 1.000 1.900 ;
        RECT  0.100 1.740 1.000 1.900 ;
        RECT  0.100 1.740 0.420 2.040 ;
        RECT  7.090 0.970 7.250 1.340 ;
        RECT  6.510 1.180 7.250 1.340 ;
        RECT  5.270 0.620 5.550 1.780 ;
        RECT  5.370 0.620 5.550 2.100 ;
        RECT  6.510 1.180 6.670 2.100 ;
        RECT  5.370 1.940 6.670 2.100 ;
        RECT  7.350 0.620 7.630 0.840 ;
        RECT  7.430 1.110 8.370 1.270 ;
        RECT  7.430 0.620 7.630 2.100 ;
        RECT  7.030 0.300 7.950 0.460 ;
        RECT  7.030 0.300 7.190 0.670 ;
        RECT  6.070 0.500 7.190 0.670 ;
        RECT  7.790 0.300 7.950 0.950 ;
        RECT  8.550 0.410 8.810 0.790 ;
        RECT  7.790 0.790 8.710 0.950 ;
        RECT  6.070 0.500 6.350 1.770 ;
        RECT  8.550 0.410 8.710 2.090 ;
        RECT  8.410 1.440 8.710 2.090 ;
        LAYER VTPH ;
        RECT  3.490 1.140 4.670 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.490 1.200 11.600 2.400 ;
        RECT  6.370 1.140 11.600 2.400 ;
        RECT  0.000 1.210 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.140 ;
        RECT  4.670 0.000 6.370 1.200 ;
        RECT  2.390 0.000 3.490 1.210 ;
    END
END DFCQM8HM

MACRO DFCQM4HM
    CLASS CORE ;
    FOREIGN DFCQM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.107  LAYER ME1  ;
        ANTENNAGATEAREA 0.107  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.378  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.240 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.564  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.030 0.830 9.560 1.160 ;
        RECT  9.030 0.390 9.230 2.100 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.580 1.410 9.740 2.540 ;
        RECT  8.370 1.420 8.570 2.540 ;
        RECT  7.370 1.460 7.570 2.540 ;
        RECT  3.780 2.000 3.980 2.540 ;
        RECT  1.780 1.750 1.980 2.540 ;
        RECT  0.660 2.060 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.550 -0.140 9.750 0.660 ;
        RECT  8.510 -0.140 8.710 0.670 ;
        RECT  7.530 -0.140 7.690 0.630 ;
        RECT  3.860 -0.140 4.140 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.120 1.120 4.400 1.340 ;
        RECT  3.060 1.290 4.280 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.620 0.620 4.910 0.950 ;
        RECT  3.640 0.800 4.720 0.960 ;
        RECT  3.640 0.800 3.920 1.100 ;
        RECT  4.560 0.800 4.720 1.780 ;
        RECT  4.500 1.500 4.780 1.780 ;
        RECT  1.340 0.620 1.620 1.570 ;
        RECT  1.340 1.400 2.300 1.570 ;
        RECT  3.440 1.680 4.340 1.840 ;
        RECT  2.140 1.400 2.300 2.090 ;
        RECT  4.180 1.680 4.340 2.100 ;
        RECT  1.340 0.620 1.500 2.080 ;
        RECT  1.260 1.720 1.500 2.080 ;
        RECT  3.440 1.680 3.600 2.090 ;
        RECT  2.140 1.930 3.600 2.090 ;
        RECT  4.180 1.940 5.190 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.580 0.460 ;
        RECT  4.300 0.300 5.910 0.460 ;
        RECT  3.400 0.300 3.580 0.640 ;
        RECT  4.300 0.300 4.460 0.640 ;
        RECT  3.400 0.480 4.460 0.640 ;
        RECT  0.140 0.300 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.750 0.300 5.910 1.700 ;
        RECT  0.800 0.750 1.000 1.900 ;
        RECT  0.100 1.740 1.000 1.900 ;
        RECT  0.100 1.740 0.420 2.040 ;
        RECT  5.270 0.620 5.550 1.780 ;
        RECT  5.370 0.620 5.550 2.100 ;
        RECT  6.510 0.970 6.670 2.100 ;
        RECT  5.370 1.940 6.670 2.100 ;
        RECT  6.770 0.620 7.050 0.840 ;
        RECT  6.850 1.110 7.810 1.270 ;
        RECT  6.850 0.620 7.050 2.100 ;
        RECT  6.070 0.300 7.370 0.460 ;
        RECT  7.210 0.300 7.370 0.950 ;
        RECT  7.970 0.490 8.270 0.790 ;
        RECT  7.210 0.790 8.130 0.950 ;
        RECT  6.070 0.300 6.350 1.770 ;
        RECT  7.970 0.490 8.130 2.090 ;
        RECT  7.830 1.440 8.130 2.090 ;
        LAYER VTPH ;
        RECT  3.490 1.140 4.670 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.490 1.200 10.000 2.400 ;
        RECT  6.370 1.140 10.000 2.400 ;
        RECT  0.000 1.210 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  4.670 0.000 6.370 1.200 ;
        RECT  2.390 0.000 3.490 1.210 ;
    END
END DFCQM4HM

MACRO DFCQM2HM
    CLASS CORE ;
    FOREIGN DFCQM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.461  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.240 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.500 0.390 8.750 1.970 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.110 1.630 9.270 2.540 ;
        RECT  7.410 1.440 7.610 2.540 ;
        RECT  3.820 2.000 4.020 2.540 ;
        RECT  1.740 1.750 1.940 2.540 ;
        RECT  0.660 2.060 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.070 -0.140 9.270 0.660 ;
        RECT  7.570 -0.140 7.730 0.630 ;
        RECT  3.900 -0.140 4.180 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.160 1.120 4.440 1.340 ;
        RECT  3.060 1.290 4.320 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.660 0.620 4.950 0.950 ;
        RECT  3.680 0.800 4.760 0.960 ;
        RECT  3.680 0.800 3.960 1.100 ;
        RECT  4.600 0.800 4.760 1.780 ;
        RECT  4.540 1.500 4.820 1.780 ;
        RECT  1.340 0.620 1.620 1.570 ;
        RECT  1.340 1.400 2.300 1.570 ;
        RECT  3.380 1.680 4.380 1.840 ;
        RECT  2.140 1.400 2.300 2.090 ;
        RECT  4.220 1.680 4.380 2.100 ;
        RECT  1.340 0.620 1.500 2.080 ;
        RECT  1.260 1.720 1.500 2.080 ;
        RECT  3.380 1.680 3.540 2.090 ;
        RECT  2.140 1.930 3.540 2.090 ;
        RECT  4.220 1.940 5.230 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.620 0.460 ;
        RECT  4.340 0.300 5.950 0.460 ;
        RECT  3.440 0.300 3.620 0.640 ;
        RECT  4.340 0.300 4.500 0.640 ;
        RECT  3.440 0.480 4.500 0.640 ;
        RECT  0.140 0.300 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.790 0.300 5.950 1.700 ;
        RECT  0.800 0.750 1.000 1.900 ;
        RECT  0.100 1.740 1.000 1.900 ;
        RECT  0.100 1.740 0.420 2.040 ;
        RECT  5.310 0.620 5.590 1.780 ;
        RECT  5.410 0.620 5.590 2.100 ;
        RECT  6.550 0.970 6.710 2.100 ;
        RECT  5.410 1.940 6.710 2.100 ;
        RECT  6.810 0.620 7.090 0.840 ;
        RECT  6.890 1.110 7.870 1.270 ;
        RECT  6.890 0.620 7.090 1.750 ;
        RECT  6.110 0.300 7.410 0.460 ;
        RECT  7.250 0.300 7.410 0.950 ;
        RECT  8.030 0.310 8.310 0.950 ;
        RECT  7.250 0.790 8.310 0.950 ;
        RECT  8.030 0.310 8.190 1.720 ;
        RECT  7.870 1.440 8.190 1.720 ;
        RECT  6.110 0.300 6.390 1.770 ;
        LAYER VTPH ;
        RECT  3.530 1.140 4.710 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.530 1.200 9.600 2.400 ;
        RECT  6.410 1.140 9.600 2.400 ;
        RECT  0.000 1.210 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  4.710 0.000 6.410 1.200 ;
        RECT  2.390 0.000 3.530 1.210 ;
    END
END DFCQM2HM

MACRO DFCQM1HM
    CLASS CORE ;
    FOREIGN DFCQM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.461  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.240 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.068  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.500 0.390 8.760 1.870 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.090 1.620 9.250 2.540 ;
        RECT  7.410 1.440 7.610 2.540 ;
        RECT  3.820 2.000 4.020 2.540 ;
        RECT  1.740 1.750 1.940 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.070 -0.140 9.270 0.660 ;
        RECT  7.570 -0.140 7.730 0.630 ;
        RECT  3.900 -0.140 4.180 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.160 1.120 4.440 1.340 ;
        RECT  3.060 1.290 4.320 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.660 0.620 4.950 0.950 ;
        RECT  3.680 0.800 4.760 0.960 ;
        RECT  3.680 0.800 3.960 1.100 ;
        RECT  4.600 0.800 4.760 1.780 ;
        RECT  4.540 1.500 4.820 1.780 ;
        RECT  1.340 0.620 1.620 1.570 ;
        RECT  1.340 1.400 2.300 1.570 ;
        RECT  3.380 1.680 4.380 1.840 ;
        RECT  2.140 1.400 2.300 2.090 ;
        RECT  4.220 1.680 4.380 2.100 ;
        RECT  1.340 0.620 1.500 2.080 ;
        RECT  1.260 1.720 1.500 2.080 ;
        RECT  3.380 1.680 3.540 2.090 ;
        RECT  2.140 1.930 3.540 2.090 ;
        RECT  4.220 1.940 5.230 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.620 0.460 ;
        RECT  4.340 0.300 5.950 0.460 ;
        RECT  3.440 0.300 3.620 0.640 ;
        RECT  4.340 0.300 4.500 0.640 ;
        RECT  3.440 0.480 4.500 0.640 ;
        RECT  0.140 0.300 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.790 0.300 5.950 1.700 ;
        RECT  0.800 0.750 1.000 1.890 ;
        RECT  0.100 1.730 1.000 1.890 ;
        RECT  0.100 1.730 0.420 2.040 ;
        RECT  5.310 0.620 5.590 1.780 ;
        RECT  5.410 0.620 5.590 2.100 ;
        RECT  6.550 0.970 6.710 2.100 ;
        RECT  5.410 1.940 6.710 2.100 ;
        RECT  6.810 0.620 7.090 0.840 ;
        RECT  6.890 1.110 7.870 1.270 ;
        RECT  6.890 0.620 7.090 1.750 ;
        RECT  6.110 0.300 7.410 0.460 ;
        RECT  8.030 0.310 8.310 0.600 ;
        RECT  7.250 0.300 7.410 0.950 ;
        RECT  7.250 0.790 8.190 0.950 ;
        RECT  8.030 0.310 8.190 1.710 ;
        RECT  7.870 1.440 8.190 1.710 ;
        RECT  6.110 0.300 6.390 1.770 ;
        LAYER VTPH ;
        RECT  3.530 1.140 4.710 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.530 1.200 9.600 2.400 ;
        RECT  6.410 1.140 9.600 2.400 ;
        RECT  0.000 1.210 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  4.710 0.000 6.410 1.200 ;
        RECT  2.390 0.000 3.530 1.210 ;
    END
END DFCQM1HM

MACRO DFCM8HM
    CLASS CORE ;
    FOREIGN DFCM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        ANTENNAGATEAREA 0.118  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.793  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.280 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.222  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.960 0.380 11.120 1.780 ;
        RECT  9.630 0.850 11.120 1.100 ;
        RECT  9.750 0.390 9.950 1.100 ;
        RECT  9.630 0.830 9.830 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  13.140 0.380 13.340 1.820 ;
        RECT  12.100 0.840 13.340 1.160 ;
        RECT  12.100 0.380 12.300 1.820 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 14.000 2.540 ;
        RECT  13.660 1.480 13.860 2.540 ;
        RECT  12.620 1.480 12.820 2.540 ;
        RECT  11.600 1.440 11.760 2.540 ;
        RECT  10.320 1.800 10.480 2.540 ;
        RECT  8.950 1.840 9.150 2.540 ;
        RECT  7.950 1.460 8.150 2.540 ;
        RECT  6.830 1.520 7.110 2.540 ;
        RECT  3.780 2.000 3.980 2.540 ;
        RECT  1.780 1.790 1.980 2.540 ;
        RECT  0.660 2.060 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 14.000 0.140 ;
        RECT  13.660 -0.140 13.860 0.660 ;
        RECT  12.620 -0.140 12.820 0.660 ;
        RECT  11.520 -0.140 11.720 0.660 ;
        RECT  10.270 -0.140 10.480 0.610 ;
        RECT  9.230 -0.140 9.430 0.610 ;
        RECT  8.110 -0.140 8.270 0.630 ;
        RECT  6.590 -0.140 6.870 0.320 ;
        RECT  3.860 -0.140 4.140 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.120 1.120 4.400 1.340 ;
        RECT  3.060 1.290 4.280 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.620 0.620 4.910 0.950 ;
        RECT  3.640 0.800 4.720 0.960 ;
        RECT  3.640 0.800 3.920 1.100 ;
        RECT  4.560 0.800 4.720 1.780 ;
        RECT  4.500 1.500 4.780 1.780 ;
        RECT  1.340 0.620 1.620 1.610 ;
        RECT  1.340 1.440 2.300 1.610 ;
        RECT  1.260 1.500 1.500 1.820 ;
        RECT  3.440 1.680 4.340 1.840 ;
        RECT  2.140 1.440 2.300 2.090 ;
        RECT  4.180 1.680 4.340 2.100 ;
        RECT  3.440 1.680 3.600 2.090 ;
        RECT  2.140 1.930 3.600 2.090 ;
        RECT  4.180 1.940 5.190 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.580 0.460 ;
        RECT  4.300 0.300 5.910 0.460 ;
        RECT  3.400 0.300 3.580 0.640 ;
        RECT  4.300 0.300 4.460 0.640 ;
        RECT  3.400 0.480 4.460 0.640 ;
        RECT  0.140 0.450 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.750 0.300 5.910 1.700 ;
        RECT  0.800 0.750 1.000 1.900 ;
        RECT  0.100 1.740 1.000 1.900 ;
        RECT  0.100 1.740 0.420 2.040 ;
        RECT  7.090 0.970 7.250 1.340 ;
        RECT  6.510 1.180 7.250 1.340 ;
        RECT  5.270 0.620 5.550 1.780 ;
        RECT  5.370 0.620 5.550 2.100 ;
        RECT  6.510 1.180 6.670 2.100 ;
        RECT  5.370 1.940 6.670 2.100 ;
        RECT  7.350 0.620 7.630 0.840 ;
        RECT  7.430 1.110 8.720 1.270 ;
        RECT  7.430 0.620 7.630 2.100 ;
        RECT  7.030 0.300 7.950 0.460 ;
        RECT  7.030 0.300 7.190 0.670 ;
        RECT  6.070 0.500 7.190 0.670 ;
        RECT  7.790 0.300 7.950 0.950 ;
        RECT  8.610 0.490 8.810 0.950 ;
        RECT  7.790 0.790 9.470 0.950 ;
        RECT  11.280 1.030 11.840 1.230 ;
        RECT  8.410 1.440 9.470 1.600 ;
        RECT  10.000 1.480 10.800 1.640 ;
        RECT  6.070 0.500 6.350 1.770 ;
        RECT  9.310 0.790 9.470 2.100 ;
        RECT  10.640 1.480 10.800 2.100 ;
        RECT  8.410 1.440 8.710 2.090 ;
        RECT  10.000 1.480 10.160 2.100 ;
        RECT  9.310 1.940 10.160 2.100 ;
        RECT  11.280 1.030 11.440 2.100 ;
        RECT  10.640 1.940 11.440 2.100 ;
        LAYER VTPH ;
        RECT  3.490 1.140 4.670 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.490 1.200 14.000 2.400 ;
        RECT  6.370 1.140 14.000 2.400 ;
        RECT  0.000 1.210 14.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 14.000 1.140 ;
        RECT  4.670 0.000 6.370 1.200 ;
        RECT  2.390 0.000 3.490 1.210 ;
    END
END DFCM8HM

MACRO DFCM4HM
    CLASS CORE ;
    FOREIGN DFCM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.107  LAYER ME1  ;
        ANTENNAGATEAREA 0.107  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.378  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.240 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.578  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.050 0.830 9.560 1.160 ;
        RECT  9.170 0.390 9.370 1.160 ;
        RECT  9.050 0.830 9.250 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.230 0.840 10.860 1.160 ;
        RECT  10.230 0.380 10.430 1.820 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.750 1.480 10.950 2.540 ;
        RECT  9.730 1.800 9.890 2.540 ;
        RECT  8.370 1.840 8.570 2.540 ;
        RECT  7.370 1.460 7.570 2.540 ;
        RECT  3.780 2.000 3.980 2.540 ;
        RECT  1.780 1.750 1.980 2.540 ;
        RECT  0.660 2.060 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.750 -0.140 10.950 0.660 ;
        RECT  9.690 -0.140 9.890 0.660 ;
        RECT  8.650 -0.140 8.850 0.610 ;
        RECT  7.530 -0.140 7.690 0.630 ;
        RECT  3.860 -0.140 4.140 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.120 1.120 4.400 1.340 ;
        RECT  3.060 1.290 4.280 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.620 0.620 4.910 0.950 ;
        RECT  3.640 0.800 4.720 0.960 ;
        RECT  3.640 0.800 3.920 1.100 ;
        RECT  4.560 0.800 4.720 1.780 ;
        RECT  4.500 1.500 4.780 1.780 ;
        RECT  1.340 0.620 1.620 1.570 ;
        RECT  1.340 1.400 2.300 1.570 ;
        RECT  3.440 1.680 4.340 1.840 ;
        RECT  2.140 1.400 2.300 2.090 ;
        RECT  4.180 1.680 4.340 2.100 ;
        RECT  1.340 0.620 1.500 2.080 ;
        RECT  1.260 1.720 1.500 2.080 ;
        RECT  3.440 1.680 3.600 2.090 ;
        RECT  2.140 1.930 3.600 2.090 ;
        RECT  4.180 1.940 5.190 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.580 0.460 ;
        RECT  4.300 0.300 5.910 0.460 ;
        RECT  3.400 0.300 3.580 0.640 ;
        RECT  4.300 0.300 4.460 0.640 ;
        RECT  3.400 0.480 4.460 0.640 ;
        RECT  0.140 0.300 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.750 0.300 5.910 1.700 ;
        RECT  0.800 0.750 1.000 1.900 ;
        RECT  0.100 1.740 1.000 1.900 ;
        RECT  0.100 1.740 0.420 2.040 ;
        RECT  5.270 0.620 5.550 1.780 ;
        RECT  5.370 0.620 5.550 2.100 ;
        RECT  6.510 0.970 6.670 2.100 ;
        RECT  5.370 1.940 6.670 2.100 ;
        RECT  6.770 0.620 7.050 0.840 ;
        RECT  6.850 1.110 8.140 1.270 ;
        RECT  6.850 0.620 7.050 2.100 ;
        RECT  6.070 0.300 7.370 0.460 ;
        RECT  7.210 0.300 7.370 0.950 ;
        RECT  8.030 0.490 8.230 0.950 ;
        RECT  7.210 0.790 8.890 0.950 ;
        RECT  7.830 1.440 8.890 1.600 ;
        RECT  9.890 0.920 10.050 1.640 ;
        RECT  9.410 1.480 10.050 1.640 ;
        RECT  6.070 0.300 6.350 1.770 ;
        RECT  8.730 0.790 8.890 2.100 ;
        RECT  7.830 1.440 8.130 2.090 ;
        RECT  9.410 1.480 9.570 2.100 ;
        RECT  8.730 1.940 9.570 2.100 ;
        LAYER VTPH ;
        RECT  3.490 1.140 4.670 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.490 1.200 11.200 2.400 ;
        RECT  6.370 1.140 11.200 2.400 ;
        RECT  0.000 1.210 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
        RECT  4.670 0.000 6.370 1.200 ;
        RECT  2.390 0.000 3.490 1.210 ;
    END
END DFCM4HM

MACRO DFCM2HM
    CLASS CORE ;
    FOREIGN DFCM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.461  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.240 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.500 0.390 8.750 1.320 ;
        RECT  8.430 1.180 8.630 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.610 0.840 9.900 1.160 ;
        RECT  9.610 0.380 9.810 1.820 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.110 1.800 9.270 2.540 ;
        RECT  7.410 1.440 7.610 2.540 ;
        RECT  3.820 2.000 4.020 2.540 ;
        RECT  1.740 1.750 1.940 2.540 ;
        RECT  0.660 2.060 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.070 -0.140 9.270 0.660 ;
        RECT  7.570 -0.140 7.730 0.630 ;
        RECT  3.900 -0.140 4.180 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.160 1.120 4.440 1.340 ;
        RECT  3.060 1.290 4.320 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.660 0.620 4.950 0.950 ;
        RECT  3.680 0.800 4.760 0.960 ;
        RECT  3.680 0.800 3.960 1.100 ;
        RECT  4.600 0.800 4.760 1.780 ;
        RECT  4.540 1.500 4.820 1.780 ;
        RECT  1.340 0.620 1.620 1.570 ;
        RECT  1.340 1.400 2.300 1.570 ;
        RECT  3.380 1.680 4.380 1.840 ;
        RECT  2.140 1.400 2.300 2.090 ;
        RECT  4.220 1.680 4.380 2.100 ;
        RECT  1.340 0.620 1.500 2.080 ;
        RECT  1.260 1.720 1.500 2.080 ;
        RECT  3.380 1.680 3.540 2.090 ;
        RECT  2.140 1.930 3.540 2.090 ;
        RECT  4.220 1.940 5.230 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.620 0.460 ;
        RECT  4.340 0.300 5.950 0.460 ;
        RECT  3.440 0.300 3.620 0.640 ;
        RECT  4.340 0.300 4.500 0.640 ;
        RECT  3.440 0.480 4.500 0.640 ;
        RECT  0.140 0.300 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.790 0.300 5.950 1.700 ;
        RECT  0.800 0.750 1.000 1.900 ;
        RECT  0.100 1.740 1.000 1.900 ;
        RECT  0.100 1.740 0.420 2.040 ;
        RECT  5.310 0.620 5.590 1.780 ;
        RECT  5.410 0.620 5.590 2.100 ;
        RECT  6.550 0.970 6.710 2.100 ;
        RECT  5.410 1.940 6.710 2.100 ;
        RECT  6.810 0.620 7.090 0.840 ;
        RECT  6.890 1.110 7.870 1.270 ;
        RECT  6.890 0.620 7.090 1.750 ;
        RECT  6.110 0.300 7.410 0.460 ;
        RECT  7.250 0.300 7.410 0.950 ;
        RECT  8.030 0.310 8.310 0.950 ;
        RECT  7.250 0.790 8.310 0.950 ;
        RECT  9.270 0.920 9.430 1.640 ;
        RECT  8.790 1.480 9.430 1.640 ;
        RECT  7.870 1.440 8.190 1.720 ;
        RECT  6.110 0.300 6.390 1.770 ;
        RECT  8.030 0.310 8.190 2.100 ;
        RECT  8.790 1.480 8.950 2.100 ;
        RECT  8.030 1.940 8.950 2.100 ;
        LAYER VTPH ;
        RECT  3.530 1.140 4.710 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.530 1.200 10.000 2.400 ;
        RECT  6.410 1.140 10.000 2.400 ;
        RECT  0.000 1.210 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  4.710 0.000 6.410 1.200 ;
        RECT  2.390 0.000 3.530 1.210 ;
    END
END DFCM2HM

MACRO DFCM1HM
    CLASS CORE ;
    FOREIGN DFCM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.072  LAYER ME1  ;
        ANTENNAGATEAREA 0.072  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 9.461  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.540 1.250 2.740 1.450 ;
        LAYER ME2 ;
        RECT  2.440 0.830 2.740 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.080 2.900 1.450 ;
        RECT  1.960 1.080 2.900 1.240 ;
        END
    END D
    PIN CKB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.068  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.070 0.480 1.560 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.500 0.390 8.760 1.100 ;
        RECT  8.430 0.900 8.630 1.780 ;
        END
    END Q
    PIN QB
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.610 0.840 9.900 1.160 ;
        RECT  9.610 0.380 9.810 1.820 ;
        END
    END QB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.110 1.620 9.270 2.540 ;
        RECT  7.410 1.440 7.610 2.540 ;
        RECT  3.820 2.000 4.020 2.540 ;
        RECT  1.740 1.750 1.940 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.070 -0.140 9.270 0.660 ;
        RECT  7.570 -0.140 7.730 0.630 ;
        RECT  3.900 -0.140 4.180 0.320 ;
        RECT  2.100 -0.140 2.300 0.600 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.940 0.680 3.220 0.900 ;
        RECT  4.160 1.120 4.440 1.340 ;
        RECT  3.060 1.290 4.320 1.450 ;
        RECT  3.060 0.680 3.220 1.770 ;
        RECT  2.530 1.610 3.220 1.770 ;
        RECT  4.660 0.620 4.950 0.950 ;
        RECT  3.680 0.800 4.760 0.960 ;
        RECT  3.680 0.800 3.960 1.100 ;
        RECT  4.600 0.800 4.760 1.780 ;
        RECT  4.540 1.500 4.820 1.780 ;
        RECT  1.340 0.620 1.620 1.570 ;
        RECT  1.340 1.400 2.300 1.570 ;
        RECT  3.380 1.680 4.380 1.840 ;
        RECT  2.140 1.400 2.300 2.090 ;
        RECT  4.220 1.680 4.380 2.100 ;
        RECT  1.340 0.620 1.500 2.080 ;
        RECT  1.260 1.720 1.500 2.080 ;
        RECT  3.380 1.680 3.540 2.090 ;
        RECT  2.140 1.930 3.540 2.090 ;
        RECT  4.220 1.940 5.230 2.100 ;
        RECT  1.020 0.300 1.940 0.460 ;
        RECT  2.460 0.300 3.620 0.460 ;
        RECT  4.340 0.300 5.950 0.460 ;
        RECT  3.440 0.300 3.620 0.640 ;
        RECT  4.340 0.300 4.500 0.640 ;
        RECT  3.440 0.480 4.500 0.640 ;
        RECT  0.140 0.300 0.340 0.910 ;
        RECT  1.780 0.300 1.940 0.920 ;
        RECT  1.020 0.300 1.180 0.910 ;
        RECT  0.140 0.750 1.180 0.910 ;
        RECT  2.460 0.300 2.620 0.920 ;
        RECT  1.780 0.760 2.620 0.920 ;
        RECT  5.790 0.300 5.950 1.700 ;
        RECT  0.800 0.750 1.000 1.890 ;
        RECT  0.100 1.730 1.000 1.890 ;
        RECT  0.100 1.730 0.420 2.040 ;
        RECT  5.310 0.620 5.590 1.780 ;
        RECT  5.410 0.620 5.590 2.100 ;
        RECT  6.550 0.970 6.710 2.100 ;
        RECT  5.410 1.940 6.710 2.100 ;
        RECT  6.810 0.620 7.090 0.840 ;
        RECT  6.890 1.110 7.870 1.270 ;
        RECT  6.890 0.620 7.090 1.750 ;
        RECT  6.110 0.300 7.410 0.460 ;
        RECT  8.030 0.310 8.310 0.600 ;
        RECT  7.250 0.300 7.410 0.950 ;
        RECT  7.250 0.790 8.190 0.950 ;
        RECT  9.270 0.920 9.430 1.420 ;
        RECT  8.790 1.260 9.430 1.420 ;
        RECT  7.870 1.440 8.190 1.720 ;
        RECT  6.110 0.300 6.390 1.770 ;
        RECT  8.030 0.310 8.190 2.100 ;
        RECT  8.790 1.260 8.950 2.100 ;
        RECT  8.030 1.940 8.950 2.100 ;
        LAYER VTPH ;
        RECT  3.530 1.140 4.710 2.400 ;
        RECT  0.000 1.140 2.390 2.400 ;
        RECT  3.530 1.200 10.000 2.400 ;
        RECT  6.410 1.140 10.000 2.400 ;
        RECT  0.000 1.210 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  4.710 0.000 6.410 1.200 ;
        RECT  2.390 0.000 3.530 1.210 ;
    END
END DFCM1HM

MACRO DEL4M4HM
    CLASS CORE ;
    FOREIGN DEL4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.097  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.660 3.900 1.500 ;
        RECT  3.500 1.300 3.700 2.100 ;
        RECT  3.500 0.330 3.700 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.720 4.220 2.540 ;
        RECT  2.980 1.530 3.180 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.610 ;
        RECT  2.980 -0.140 3.180 0.610 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.360 0.680 ;
        RECT  1.200 0.520 1.360 1.480 ;
        RECT  0.160 1.320 1.360 1.480 ;
        RECT  0.160 1.320 0.320 1.850 ;
        RECT  1.640 0.360 1.820 1.140 ;
        RECT  1.640 0.930 2.460 1.140 ;
        RECT  1.640 0.360 1.800 1.850 ;
        RECT  2.020 0.420 2.820 0.580 ;
        RECT  2.620 0.980 3.540 1.140 ;
        RECT  2.620 0.420 2.820 1.750 ;
        RECT  2.020 1.590 2.820 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END DEL4M4HM

MACRO DEL4M1HM
    CLASS CORE ;
    FOREIGN DEL4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.046  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.281  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.560 3.900 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.060 1.940 3.260 2.540 ;
        RECT  0.700 1.640 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.260 0.400 ;
        RECT  0.700 -0.140 0.980 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.400 0.680 ;
        RECT  1.240 0.520 1.400 1.480 ;
        RECT  0.160 1.320 1.400 1.480 ;
        RECT  0.160 1.320 0.320 1.900 ;
        RECT  1.720 1.060 2.940 1.220 ;
        RECT  1.720 0.340 1.880 1.900 ;
        RECT  2.100 0.620 3.460 0.780 ;
        RECT  3.300 0.620 3.460 1.660 ;
        RECT  2.100 1.500 3.460 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END DEL4M1HM

MACRO DEL3M4HM
    CLASS CORE ;
    FOREIGN DEL3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.097  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.660 3.900 1.500 ;
        RECT  3.500 1.300 3.700 2.100 ;
        RECT  3.500 0.330 3.700 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.720 4.220 2.540 ;
        RECT  2.980 1.530 3.180 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.610 ;
        RECT  2.980 -0.140 3.180 0.610 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.360 0.680 ;
        RECT  1.200 0.520 1.360 1.480 ;
        RECT  0.160 1.320 1.360 1.480 ;
        RECT  0.160 1.320 0.320 1.850 ;
        RECT  1.640 0.360 1.820 1.140 ;
        RECT  1.640 0.930 2.460 1.140 ;
        RECT  1.640 0.360 1.800 1.850 ;
        RECT  2.020 0.420 2.820 0.580 ;
        RECT  2.620 0.980 3.540 1.140 ;
        RECT  2.620 0.420 2.820 1.750 ;
        RECT  2.020 1.590 2.820 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END DEL3M4HM

MACRO DEL3M1HM
    CLASS CORE ;
    FOREIGN DEL3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.046  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.281  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.560 3.900 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.060 1.940 3.260 2.540 ;
        RECT  0.700 1.640 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.260 0.400 ;
        RECT  0.700 -0.140 0.980 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.400 0.680 ;
        RECT  1.240 0.520 1.400 1.480 ;
        RECT  0.160 1.320 1.400 1.480 ;
        RECT  0.160 1.320 0.320 1.900 ;
        RECT  1.720 1.060 2.940 1.220 ;
        RECT  1.720 0.340 1.880 1.900 ;
        RECT  2.100 0.620 3.460 0.780 ;
        RECT  3.300 0.620 3.460 1.660 ;
        RECT  2.100 1.500 3.460 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END DEL3M1HM

MACRO DEL2M4HM
    CLASS CORE ;
    FOREIGN DEL2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.097  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.660 3.900 1.500 ;
        RECT  3.500 1.300 3.700 2.100 ;
        RECT  3.500 0.330 3.700 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.720 4.220 2.540 ;
        RECT  2.980 1.530 3.180 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.610 ;
        RECT  2.980 -0.140 3.180 0.610 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.360 0.680 ;
        RECT  1.200 0.520 1.360 1.480 ;
        RECT  0.160 1.320 1.360 1.480 ;
        RECT  0.160 1.320 0.320 1.850 ;
        RECT  1.640 0.360 1.820 1.140 ;
        RECT  1.640 0.930 2.460 1.140 ;
        RECT  1.640 0.360 1.800 1.850 ;
        RECT  2.020 0.420 2.820 0.580 ;
        RECT  2.620 0.980 3.540 1.140 ;
        RECT  2.620 0.420 2.820 1.750 ;
        RECT  2.020 1.590 2.820 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END DEL2M4HM

MACRO DEL2M1HM
    CLASS CORE ;
    FOREIGN DEL2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.046  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.281  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.560 3.900 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.060 1.940 3.260 2.540 ;
        RECT  0.700 1.640 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.260 0.400 ;
        RECT  0.700 -0.140 0.980 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.400 0.680 ;
        RECT  1.240 0.520 1.400 1.480 ;
        RECT  0.160 1.320 1.400 1.480 ;
        RECT  0.160 1.320 0.320 1.900 ;
        RECT  1.720 1.060 2.940 1.220 ;
        RECT  1.720 0.340 1.880 1.900 ;
        RECT  2.100 0.620 3.460 0.780 ;
        RECT  3.300 0.620 3.460 1.660 ;
        RECT  2.100 1.500 3.460 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END DEL2M1HM

MACRO DEL1M4HM
    CLASS CORE ;
    FOREIGN DEL1M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.097  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.700 0.660 3.900 1.500 ;
        RECT  3.500 1.300 3.700 2.100 ;
        RECT  3.500 0.330 3.700 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.020 1.720 4.220 2.540 ;
        RECT  2.980 1.530 3.180 2.540 ;
        RECT  0.660 1.640 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.610 ;
        RECT  2.980 -0.140 3.180 0.610 ;
        RECT  0.660 -0.140 0.940 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.360 0.680 ;
        RECT  1.200 0.520 1.360 1.480 ;
        RECT  0.160 1.320 1.360 1.480 ;
        RECT  0.160 1.320 0.320 1.850 ;
        RECT  1.640 0.360 1.820 1.140 ;
        RECT  1.640 0.930 2.460 1.140 ;
        RECT  1.640 0.360 1.800 1.850 ;
        RECT  2.020 0.420 2.820 0.580 ;
        RECT  2.620 0.980 3.540 1.140 ;
        RECT  2.620 0.420 2.820 1.750 ;
        RECT  2.020 1.590 2.820 1.750 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END DEL1M4HM

MACRO DEL1M1HM
    CLASS CORE ;
    FOREIGN DEL1M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.046  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.380 0.840 0.700 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.281  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.560 3.900 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.060 1.940 3.260 2.540 ;
        RECT  0.700 1.640 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.060 -0.140 3.260 0.400 ;
        RECT  0.700 -0.140 0.980 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.320 0.320 0.680 ;
        RECT  0.160 0.520 1.400 0.680 ;
        RECT  1.240 0.520 1.400 1.480 ;
        RECT  0.160 1.320 1.400 1.480 ;
        RECT  0.160 1.320 0.320 1.900 ;
        RECT  1.720 1.060 2.940 1.220 ;
        RECT  1.720 0.340 1.880 1.900 ;
        RECT  2.100 0.620 3.460 0.780 ;
        RECT  3.300 0.620 3.460 1.660 ;
        RECT  2.100 1.500 3.460 1.660 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END DEL1M1HM

MACRO CKXOR2M8HM
    CLASS CORE ;
    FOREIGN CKXOR2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        ANTENNAGATEAREA 0.220  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.752  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.120 1.020 4.320 1.220 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.320 1.540 ;
        LAYER ME1 ;
        RECT  4.120 0.880 4.380 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.228  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 1.100 1.280 ;
        RECT  0.100 0.840 0.300 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.825  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.940 1.450 6.300 2.030 ;
        RECT  6.100 0.360 6.300 2.030 ;
        RECT  4.900 0.680 6.300 0.880 ;
        RECT  5.940 0.360 6.300 0.880 ;
        RECT  4.860 1.450 6.300 1.650 ;
        RECT  4.900 0.360 5.100 0.880 ;
        RECT  4.860 1.450 5.080 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.460 1.780 6.660 2.540 ;
        RECT  5.380 1.810 5.660 2.540 ;
        RECT  4.400 1.840 4.600 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.720 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.380 -0.140 5.660 0.520 ;
        RECT  4.380 -0.140 4.580 0.680 ;
        RECT  1.160 -0.140 1.360 0.580 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.840 0.620 2.120 0.930 ;
        RECT  1.840 0.620 2.000 2.060 ;
        RECT  1.620 1.900 2.000 2.060 ;
        RECT  1.520 0.300 2.980 0.460 ;
        RECT  0.640 0.310 0.870 0.900 ;
        RECT  2.810 0.600 3.170 0.890 ;
        RECT  1.520 0.300 1.680 0.900 ;
        RECT  0.640 0.740 1.680 0.900 ;
        RECT  2.810 0.300 2.980 1.780 ;
        RECT  1.380 0.740 1.540 1.740 ;
        RECT  0.580 1.580 1.540 1.740 ;
        RECT  2.700 1.560 3.060 1.780 ;
        RECT  3.760 0.470 4.140 0.630 ;
        RECT  3.150 1.110 3.920 1.390 ;
        RECT  3.760 0.470 3.920 1.690 ;
        RECT  2.300 0.620 2.650 0.890 ;
        RECT  4.540 1.080 5.920 1.280 ;
        RECT  4.540 1.080 4.700 1.680 ;
        RECT  4.080 1.520 4.700 1.680 ;
        RECT  2.300 0.620 2.490 2.100 ;
        RECT  2.240 1.730 2.490 2.100 ;
        RECT  3.340 1.770 3.540 2.100 ;
        RECT  4.080 1.520 4.240 2.100 ;
        RECT  2.240 1.940 4.240 2.100 ;
        LAYER VTPH ;
        RECT  3.470 1.010 4.460 2.400 ;
        RECT  3.380 1.110 4.460 2.400 ;
        RECT  0.000 1.140 1.500 2.400 ;
        RECT  3.380 1.140 6.800 2.400 ;
        RECT  0.000 1.190 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.010 ;
        RECT  0.000 0.000 3.470 1.110 ;
        RECT  0.000 0.000 3.380 1.140 ;
        RECT  4.460 0.000 6.800 1.140 ;
        RECT  1.500 0.000 3.380 1.190 ;
    END
END CKXOR2M8HM

MACRO CKXOR2M4HM
    CLASS CORE ;
    FOREIGN CKXOR2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.120  LAYER ME1  ;
        ANTENNAGATEAREA 0.120  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.553  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.490 0.950 0.700 1.600 ;
        LAYER ME1 ;
        RECT  0.200 1.080 0.700 1.400 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.640 0.760 3.940 1.340 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.400  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.420 1.540 5.100 1.740 ;
        RECT  4.900 0.700 5.100 1.740 ;
        RECT  4.460 0.700 5.100 0.900 ;
        RECT  4.460 0.330 4.660 0.900 ;
        RECT  4.420 1.540 4.640 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  4.940 1.900 5.220 2.540 ;
        RECT  3.960 1.840 4.160 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  4.940 -0.140 5.220 0.540 ;
        RECT  3.940 -0.140 4.140 0.600 ;
        RECT  0.640 -0.140 0.840 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.600 0.880 ;
        RECT  1.320 0.620 1.480 2.050 ;
        RECT  1.100 1.890 1.480 2.050 ;
        RECT  1.000 0.300 2.460 0.460 ;
        RECT  2.290 0.300 2.460 0.840 ;
        RECT  0.160 0.300 0.320 0.900 ;
        RECT  2.290 0.640 2.640 0.840 ;
        RECT  1.000 0.300 1.160 0.900 ;
        RECT  0.160 0.740 1.160 0.900 ;
        RECT  2.290 0.300 2.450 1.780 ;
        RECT  0.860 0.740 1.020 1.740 ;
        RECT  0.100 1.580 1.020 1.740 ;
        RECT  2.160 1.540 2.540 1.780 ;
        RECT  0.100 1.580 0.320 1.990 ;
        RECT  3.320 0.380 3.700 0.540 ;
        RECT  2.670 1.100 3.480 1.380 ;
        RECT  3.320 0.380 3.480 1.760 ;
        RECT  1.760 0.620 2.130 0.880 ;
        RECT  4.100 1.080 4.710 1.280 ;
        RECT  4.100 1.080 4.260 1.660 ;
        RECT  3.640 1.500 4.260 1.660 ;
        RECT  1.760 0.620 1.920 2.100 ;
        RECT  1.720 1.730 1.920 2.100 ;
        RECT  2.820 1.800 3.020 2.100 ;
        RECT  3.640 1.500 3.800 2.100 ;
        RECT  1.720 1.940 3.800 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.950 2.400 ;
        RECT  2.800 1.140 5.600 2.400 ;
        RECT  0.000 1.180 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
        RECT  0.950 0.000 2.800 1.180 ;
    END
END CKXOR2M4HM

MACRO CKXOR2M2HM
    CLASS CORE ;
    FOREIGN CKXOR2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.337  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.330 3.900 1.970 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.197  LAYER ME1  ;
        ANTENNAGATEAREA 0.197  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.982  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.060 0.700 1.260 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.420 0.970 0.820 1.320 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.780 3.160 1.350 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.160 1.830 3.400 2.540 ;
        RECT  0.640 1.800 0.880 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.140 -0.140 3.340 0.600 ;
        RECT  0.680 -0.140 0.880 0.810 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.360 0.620 1.660 0.820 ;
        RECT  1.360 0.620 1.520 1.780 ;
        RECT  0.100 0.530 0.380 0.800 ;
        RECT  1.680 1.020 1.960 1.220 ;
        RECT  0.100 0.530 0.260 1.910 ;
        RECT  0.100 1.480 1.200 1.640 ;
        RECT  0.100 1.480 0.320 1.910 ;
        RECT  1.040 1.480 1.200 2.100 ;
        RECT  1.680 1.020 1.840 2.100 ;
        RECT  1.040 1.940 1.840 2.100 ;
        RECT  1.040 0.300 2.860 0.460 ;
        RECT  2.520 0.300 2.860 0.570 ;
        RECT  1.040 0.300 1.200 1.300 ;
        RECT  2.520 0.300 2.680 1.780 ;
        RECT  1.980 0.620 2.360 0.820 ;
        RECT  3.340 0.990 3.500 1.670 ;
        RECT  2.840 1.510 3.500 1.670 ;
        RECT  2.000 1.590 2.360 1.870 ;
        RECT  2.190 0.620 2.360 2.100 ;
        RECT  2.840 1.510 3.000 2.100 ;
        RECT  2.190 1.940 3.000 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END CKXOR2M2HM

MACRO CKXOR2M1HM
    CLASS CORE ;
    FOREIGN CKXOR2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER ME1  ;
        ANTENNAGATEAREA 0.194  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.033  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.060 0.700 1.260 ;
        LAYER ME2 ;
        RECT  0.500 0.890 0.700 1.690 ;
        LAYER ME1 ;
        RECT  0.420 0.960 0.820 1.320 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.820 3.160 1.360 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.258  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.320 3.900 2.070 ;
        RECT  3.530 0.320 3.900 0.690 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.160 1.840 3.400 2.540 ;
        RECT  0.580 1.800 0.840 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.020 -0.140 3.220 0.600 ;
        RECT  0.620 -0.140 0.840 0.800 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.320 0.620 1.520 1.780 ;
        RECT  0.100 0.520 0.360 0.800 ;
        RECT  1.680 1.060 1.960 1.260 ;
        RECT  0.100 0.520 0.260 1.910 ;
        RECT  0.100 1.480 1.160 1.640 ;
        RECT  0.100 1.480 0.320 1.910 ;
        RECT  1.000 1.480 1.160 2.100 ;
        RECT  1.680 1.060 1.840 2.100 ;
        RECT  1.000 1.940 1.840 2.100 ;
        RECT  1.000 0.300 2.800 0.460 ;
        RECT  2.520 0.300 2.800 0.620 ;
        RECT  1.000 0.300 1.160 1.300 ;
        RECT  2.520 0.300 2.680 1.780 ;
        RECT  1.890 0.620 2.350 0.830 ;
        RECT  3.340 0.990 3.500 1.680 ;
        RECT  2.840 1.520 3.500 1.680 ;
        RECT  2.000 1.590 2.350 1.870 ;
        RECT  2.190 0.620 2.350 2.100 ;
        RECT  2.840 1.520 3.000 2.100 ;
        RECT  2.190 1.940 3.000 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.080 2.400 ;
        RECT  1.760 1.140 4.000 2.400 ;
        RECT  0.000 1.200 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  1.080 0.000 1.760 1.200 ;
    END
END CKXOR2M1HM

MACRO CKXOR2M12HM
    CLASS CORE ;
    FOREIGN CKXOR2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.364  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.840 6.740 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.350  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.020 1.520 1.220 ;
        RECT  0.500 0.840 0.700 1.220 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.204  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.460 1.360 9.660 2.100 ;
        RECT  7.400 0.660 9.660 0.860 ;
        RECT  9.460 0.310 9.660 0.860 ;
        RECT  7.380 1.360 9.660 1.560 ;
        RECT  8.450 0.660 8.750 1.560 ;
        RECT  8.420 1.360 8.620 2.100 ;
        RECT  8.420 0.310 8.620 0.860 ;
        RECT  7.400 0.310 7.600 0.860 ;
        RECT  7.380 1.360 7.580 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  9.980 1.720 10.180 2.540 ;
        RECT  8.940 1.720 9.140 2.540 ;
        RECT  7.900 1.720 8.100 2.540 ;
        RECT  6.860 1.720 7.060 2.540 ;
        RECT  5.780 1.860 6.060 2.540 ;
        RECT  2.820 2.080 3.100 2.540 ;
        RECT  1.700 2.080 1.980 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  8.900 -0.140 9.190 0.500 ;
        RECT  7.860 -0.140 8.140 0.500 ;
        RECT  6.780 -0.140 7.060 0.360 ;
        RECT  1.660 -0.140 1.940 0.510 ;
        RECT  0.660 -0.140 0.860 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.240 0.400 2.460 0.690 ;
        RECT  2.240 0.530 3.960 0.690 ;
        RECT  2.220 1.440 3.960 1.600 ;
        RECT  3.800 0.530 3.960 1.780 ;
        RECT  1.200 0.330 1.360 0.830 ;
        RECT  1.200 0.670 2.060 0.830 ;
        RECT  4.700 0.620 5.000 0.840 ;
        RECT  1.900 1.010 2.720 1.170 ;
        RECT  0.140 1.380 2.060 1.540 ;
        RECT  1.180 1.380 2.060 1.580 ;
        RECT  1.900 0.670 2.060 1.920 ;
        RECT  1.900 1.760 3.490 1.920 ;
        RECT  3.330 1.760 3.490 2.100 ;
        RECT  0.140 1.380 0.340 2.100 ;
        RECT  1.180 1.380 1.380 2.100 ;
        RECT  4.840 0.620 5.000 2.100 ;
        RECT  3.330 1.940 5.000 2.100 ;
        RECT  5.680 0.620 6.300 0.820 ;
        RECT  5.680 0.620 5.840 1.700 ;
        RECT  5.680 1.540 6.520 1.700 ;
        RECT  6.360 1.540 6.520 1.990 ;
        RECT  4.160 0.300 6.620 0.460 ;
        RECT  6.460 0.300 6.620 0.680 ;
        RECT  6.460 0.520 7.100 0.680 ;
        RECT  6.940 0.520 7.100 1.200 ;
        RECT  6.940 1.040 7.940 1.200 ;
        RECT  4.160 0.300 4.320 1.780 ;
        RECT  4.160 1.620 4.580 1.780 ;
        RECT  5.360 0.300 5.520 1.990 ;
        RECT  9.200 1.040 9.920 1.200 ;
        LAYER VTPH ;
        RECT  1.450 1.080 3.400 2.400 ;
        RECT  0.000 1.140 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.080 ;
        RECT  0.000 0.000 1.450 1.140 ;
        RECT  3.400 0.000 10.400 1.140 ;
    END
END CKXOR2M12HM

MACRO CKND2M8HM
    CLASS CORE ;
    FOREIGN CKND2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.563  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.250 3.880 1.410 ;
        RECT  3.600 1.120 3.880 1.410 ;
        RECT  1.520 1.120 2.160 1.410 ;
        RECT  0.500 0.840 0.700 1.410 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.563  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 0.800 4.340 1.360 ;
        RECT  1.020 0.800 4.340 0.960 ;
        RECT  2.360 0.800 3.080 1.090 ;
        RECT  1.020 0.800 1.300 1.090 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.482  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.620 1.570 4.700 1.730 ;
        RECT  4.500 0.480 4.700 1.730 ;
        RECT  1.660 0.480 4.700 0.640 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.340 -0.140 4.620 0.320 ;
        RECT  2.580 -0.140 2.860 0.320 ;
        RECT  0.900 -0.140 1.100 0.620 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  3.260 1.900 3.540 2.540 ;
        RECT  2.220 1.900 2.500 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.140 1.640 0.420 2.540 ;
        END
    END VDD
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END CKND2M8HM

MACRO CKND2M6HM
    CLASS CORE ;
    FOREIGN CKND2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.800 2.640 1.080 ;
        RECT  0.500 0.800 2.640 0.960 ;
        RECT  0.500 0.800 0.700 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.060 1.260 3.130 1.420 ;
        RECT  2.880 0.840 3.130 1.420 ;
        RECT  1.060 1.120 1.700 1.420 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.190  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.580 1.580 3.500 1.740 ;
        RECT  3.300 0.480 3.500 1.740 ;
        RECT  0.260 0.480 3.500 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  1.240 -0.140 1.520 0.320 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END CKND2M6HM

MACRO CKND2M4HM
    CLASS CORE ;
    FOREIGN CKND2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.282  LAYER ME1  ;
        ANTENNAGATEAREA 0.282  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.826  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.100 1.100 1.300 ;
        LAYER ME2 ;
        RECT  0.900 0.910 1.100 1.690 ;
        LAYER ME1 ;
        RECT  0.860 1.010 1.500 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.282  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.090 2.280 1.290 ;
        RECT  1.660 0.660 1.860 1.290 ;
        RECT  0.500 0.660 1.860 0.840 ;
        RECT  0.280 1.090 0.700 1.290 ;
        RECT  0.500 0.660 0.700 1.290 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.940  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.620 1.540 2.700 1.740 ;
        RECT  2.500 0.770 2.700 1.740 ;
        RECT  2.020 0.770 2.700 0.930 ;
        RECT  2.020 0.340 2.180 0.930 ;
        RECT  0.900 0.340 2.180 0.500 ;
        RECT  1.640 1.540 1.940 2.080 ;
        RECT  0.620 1.540 0.910 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.340 -0.140 2.580 0.610 ;
        RECT  0.140 -0.140 0.340 0.700 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END CKND2M4HM

MACRO CKND2M2HM
    CLASS CORE ;
    FOREIGN CKND2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.780 1.100 1.380 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.320 0.840 0.700 1.360 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.458  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.540 1.500 1.740 ;
        RECT  1.300 0.300 1.500 1.740 ;
        RECT  1.020 0.300 1.500 0.570 ;
        RECT  0.660 1.540 0.930 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.140 1.540 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.180 -0.140 0.380 0.590 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END CKND2M2HM

MACRO CKND2M16HM
    CLASS CORE ;
    FOREIGN CKND2M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.126  LAYER ME2  ;
        ANTENNAGATEAREA 1.126  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 3.825  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.130 3.900 1.330 ;
        LAYER ME2 ;
        RECT  3.700 0.840 3.900 1.560 ;
        LAYER ME1 ;
        RECT  0.400 1.260 7.770 1.420 ;
        RECT  7.000 1.120 7.770 1.420 ;
        RECT  2.080 1.250 7.770 1.420 ;
        RECT  5.640 1.120 5.920 1.420 ;
        RECT  3.480 1.120 4.200 1.420 ;
        RECT  2.080 1.120 2.360 1.420 ;
        RECT  0.400 1.040 0.680 1.420 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.100 0.800 8.300 1.250 ;
        RECT  0.970 0.800 8.300 0.960 ;
        RECT  6.160 0.800 6.800 1.090 ;
        RECT  4.400 0.800 5.040 1.090 ;
        RECT  3.000 0.800 3.280 1.090 ;
        RECT  0.970 0.800 1.430 1.100 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.124  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.580 1.580 8.700 1.740 ;
        RECT  8.500 0.480 8.700 1.740 ;
        RECT  0.960 0.480 8.700 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.580 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.220 -0.140 7.500 0.320 ;
        RECT  5.460 -0.140 5.740 0.320 ;
        RECT  3.700 -0.140 3.980 0.320 ;
        RECT  1.940 -0.140 2.220 0.320 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END CKND2M16HM

MACRO CKND2M12HM
    CLASS CORE ;
    FOREIGN CKND2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.790  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 0.800 6.340 1.300 ;
        RECT  0.960 0.800 6.340 0.960 ;
        RECT  4.660 0.800 4.940 1.100 ;
        RECT  2.960 0.800 3.240 1.100 ;
        RECT  0.960 0.800 1.600 1.090 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.790  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.260 5.920 1.420 ;
        RECT  5.640 1.120 5.920 1.420 ;
        RECT  3.480 1.120 4.120 1.420 ;
        RECT  2.060 1.120 2.340 1.420 ;
        RECT  0.500 0.840 0.700 1.420 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.202  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.580 6.700 1.740 ;
        RECT  6.500 0.480 6.700 1.740 ;
        RECT  2.740 0.480 6.700 0.640 ;
        RECT  5.860 1.580 6.060 1.910 ;
        RECT  4.820 1.580 5.020 1.910 ;
        RECT  3.780 1.580 3.980 1.910 ;
        RECT  2.740 1.580 2.940 1.910 ;
        RECT  1.700 1.580 1.900 1.910 ;
        RECT  0.660 1.580 0.860 1.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.420 -0.140 5.700 0.320 ;
        RECT  3.660 -0.140 3.940 0.320 ;
        RECT  1.980 -0.140 2.180 0.640 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END CKND2M12HM

MACRO CKMUX2M8HM
    CLASS CORE ;
    FOREIGN CKMUX2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.010 3.560 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.160 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.300 2.060 1.090 ;
        RECT  1.100 0.300 2.060 0.460 ;
        RECT  0.500 0.540 1.270 0.700 ;
        RECT  1.100 0.300 1.270 0.700 ;
        RECT  0.500 0.540 0.700 1.320 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.846  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.580 0.720 5.820 0.920 ;
        RECT  5.620 0.300 5.820 0.920 ;
        RECT  5.060 1.440 5.340 2.080 ;
        RECT  4.900 0.720 5.100 1.640 ;
        RECT  4.060 1.440 5.340 1.640 ;
        RECT  4.580 0.390 4.780 0.920 ;
        RECT  4.060 1.440 4.260 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.620 1.480 5.820 2.540 ;
        RECT  4.580 1.840 4.780 2.540 ;
        RECT  3.540 1.840 3.740 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.300 0.560 ;
        RECT  4.060 -0.140 4.260 0.620 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.620 1.740 0.840 ;
        RECT  1.460 0.620 1.660 1.720 ;
        RECT  0.140 0.540 0.340 1.920 ;
        RECT  0.140 1.760 1.300 1.920 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  2.540 0.710 2.700 2.100 ;
        RECT  1.140 1.940 2.700 2.100 ;
        RECT  2.860 0.620 3.140 0.840 ;
        RECT  2.860 0.620 3.020 1.930 ;
        RECT  2.860 1.730 3.260 1.930 ;
        RECT  2.220 0.300 3.900 0.460 ;
        RECT  3.720 0.300 3.900 1.280 ;
        RECT  3.720 1.080 4.520 1.280 ;
        RECT  2.220 0.300 2.380 1.720 ;
        RECT  1.940 1.560 2.380 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END CKMUX2M8HM

MACRO CKMUX2M6HM
    CLASS CORE ;
    FOREIGN CKMUX2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.010 3.560 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.160 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.300 2.060 1.090 ;
        RECT  1.100 0.300 2.060 0.460 ;
        RECT  0.500 0.540 1.270 0.700 ;
        RECT  1.100 0.300 1.270 0.700 ;
        RECT  0.500 0.540 0.700 1.320 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.697  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.100 0.720 5.300 2.080 ;
        RECT  4.060 1.440 5.300 1.640 ;
        RECT  4.840 0.720 5.300 1.640 ;
        RECT  4.580 0.720 5.300 0.920 ;
        RECT  4.580 0.390 4.780 0.920 ;
        RECT  4.060 1.440 4.260 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  4.580 1.840 4.780 2.540 ;
        RECT  3.540 1.840 3.740 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.100 -0.140 5.300 0.560 ;
        RECT  4.060 -0.140 4.260 0.620 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.620 1.740 0.840 ;
        RECT  1.460 0.620 1.660 1.720 ;
        RECT  0.140 0.540 0.340 1.920 ;
        RECT  0.140 1.760 1.300 1.920 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  2.540 0.710 2.700 2.100 ;
        RECT  1.140 1.940 2.700 2.100 ;
        RECT  2.860 0.620 3.140 0.840 ;
        RECT  2.860 0.620 3.020 1.930 ;
        RECT  2.860 1.730 3.260 1.930 ;
        RECT  2.220 0.300 3.900 0.460 ;
        RECT  3.720 0.300 3.900 1.280 ;
        RECT  3.720 1.080 4.520 1.280 ;
        RECT  2.220 0.300 2.380 1.720 ;
        RECT  1.940 1.560 2.380 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END CKMUX2M6HM

MACRO CKMUX2M4HM
    CLASS CORE ;
    FOREIGN CKMUX2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.560 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.160 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.300 2.060 1.090 ;
        RECT  1.100 0.300 2.060 0.460 ;
        RECT  0.500 0.540 1.270 0.700 ;
        RECT  1.100 0.300 1.270 0.700 ;
        RECT  0.500 0.540 0.700 1.320 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.402  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.440 4.560 1.640 ;
        RECT  4.360 0.700 4.560 1.640 ;
        RECT  4.140 0.700 4.560 0.900 ;
        RECT  4.100 1.440 4.340 2.080 ;
        RECT  4.140 0.300 4.340 0.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.660 1.840 4.860 2.540 ;
        RECT  3.580 1.840 3.780 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.660 -0.140 4.860 0.560 ;
        RECT  3.620 -0.140 3.820 0.560 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.620 1.740 0.840 ;
        RECT  1.460 0.620 1.660 1.720 ;
        RECT  0.140 0.540 0.340 1.920 ;
        RECT  0.140 1.760 1.300 1.920 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  2.540 0.710 2.700 2.100 ;
        RECT  1.140 1.940 2.700 2.100 ;
        RECT  2.860 0.620 3.140 0.840 ;
        RECT  2.860 0.620 3.020 1.930 ;
        RECT  2.860 1.730 3.260 1.930 ;
        RECT  2.220 0.300 3.460 0.460 ;
        RECT  3.300 0.300 3.460 0.880 ;
        RECT  3.300 0.720 3.880 0.880 ;
        RECT  3.720 0.720 3.880 1.280 ;
        RECT  3.720 1.080 4.200 1.280 ;
        RECT  2.220 0.300 2.380 1.720 ;
        RECT  1.940 1.560 2.380 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END CKMUX2M4HM

MACRO CKMUX2M3HM
    CLASS CORE ;
    FOREIGN CKMUX2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.560 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.160 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.300 2.060 1.090 ;
        RECT  1.100 0.300 2.060 0.460 ;
        RECT  0.500 0.540 1.270 0.700 ;
        RECT  1.100 0.300 1.270 0.700 ;
        RECT  0.500 0.540 0.700 1.320 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.373  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.440 4.560 1.640 ;
        RECT  4.360 0.420 4.560 1.640 ;
        RECT  4.100 0.420 4.560 0.620 ;
        RECT  4.100 1.440 4.340 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.660 1.840 4.860 2.540 ;
        RECT  3.580 1.840 3.780 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  3.620 -0.140 3.820 0.560 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.620 1.740 0.840 ;
        RECT  1.460 0.620 1.660 1.720 ;
        RECT  0.140 0.540 0.340 1.920 ;
        RECT  0.140 1.760 1.300 1.920 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  2.540 0.710 2.700 2.100 ;
        RECT  1.140 1.940 2.700 2.100 ;
        RECT  2.860 0.620 3.140 0.840 ;
        RECT  2.860 0.620 3.020 1.930 ;
        RECT  2.860 1.730 3.260 1.930 ;
        RECT  2.220 0.300 3.460 0.460 ;
        RECT  3.300 0.300 3.460 0.880 ;
        RECT  3.300 0.720 3.880 0.880 ;
        RECT  3.720 0.720 3.880 1.280 ;
        RECT  3.720 1.080 4.200 1.280 ;
        RECT  2.220 0.300 2.380 1.720 ;
        RECT  1.940 1.560 2.380 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END CKMUX2M3HM

MACRO CKMUX2M2HM
    CLASS CORE ;
    FOREIGN CKMUX2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.560 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.160 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.300 2.060 1.090 ;
        RECT  1.100 0.300 2.060 0.460 ;
        RECT  0.500 0.540 1.270 0.700 ;
        RECT  1.100 0.300 1.270 0.700 ;
        RECT  0.500 0.540 0.700 1.320 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.340  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.520 4.400 2.100 ;
        RECT  4.200 0.360 4.400 2.100 ;
        RECT  4.100 0.360 4.400 0.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.580 1.840 3.780 2.540 ;
        RECT  0.700 2.080 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.620 -0.140 3.820 0.560 ;
        RECT  0.740 -0.140 0.940 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.460 0.620 1.740 0.840 ;
        RECT  1.460 0.620 1.660 1.780 ;
        RECT  0.140 0.540 0.340 1.920 ;
        RECT  0.140 1.760 1.300 1.920 ;
        RECT  1.140 1.760 1.300 2.100 ;
        RECT  2.540 0.710 2.700 2.100 ;
        RECT  1.140 1.940 2.700 2.100 ;
        RECT  2.860 0.620 3.140 0.840 ;
        RECT  2.860 0.620 3.020 1.930 ;
        RECT  2.860 1.730 3.260 1.930 ;
        RECT  2.220 0.300 3.460 0.460 ;
        RECT  3.300 0.300 3.460 0.880 ;
        RECT  3.300 0.720 4.040 0.880 ;
        RECT  3.840 0.720 4.040 1.180 ;
        RECT  2.220 0.300 2.380 1.720 ;
        RECT  1.940 1.560 2.380 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END CKMUX2M2HM

MACRO CKMUX2M12HM
    CLASS CORE ;
    FOREIGN CKMUX2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.114  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.120 1.050 3.500 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.109  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.080 1.140 1.560 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.161  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.740 0.320 1.900 1.090 ;
        RECT  0.970 0.320 1.900 0.480 ;
        RECT  0.500 0.540 1.140 0.700 ;
        RECT  0.970 0.320 1.140 0.700 ;
        RECT  0.500 0.540 0.700 1.320 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.164  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.930 1.440 6.140 2.080 ;
        RECT  4.900 0.720 6.140 0.920 ;
        RECT  5.940 0.390 6.140 0.920 ;
        RECT  3.860 1.440 6.140 1.640 ;
        RECT  5.660 0.720 5.900 1.640 ;
        RECT  4.900 1.440 5.100 2.080 ;
        RECT  4.900 0.390 5.100 0.920 ;
        RECT  3.860 1.440 4.060 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.460 1.480 6.660 2.540 ;
        RECT  5.420 1.840 5.620 2.540 ;
        RECT  4.380 1.840 4.580 2.540 ;
        RECT  3.340 1.840 3.540 2.540 ;
        RECT  0.530 2.080 0.810 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.460 -0.140 6.660 0.670 ;
        RECT  5.420 -0.140 5.620 0.560 ;
        RECT  4.380 -0.140 4.580 0.620 ;
        RECT  4.020 -0.140 4.220 0.620 ;
        RECT  0.610 -0.140 0.810 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.300 0.640 1.580 0.860 ;
        RECT  1.300 0.640 1.500 1.740 ;
        RECT  0.140 0.540 0.340 1.920 ;
        RECT  0.140 1.760 1.130 1.920 ;
        RECT  2.380 0.710 2.540 2.080 ;
        RECT  0.970 1.920 2.540 2.080 ;
        RECT  2.700 0.640 2.980 0.860 ;
        RECT  2.700 0.640 2.860 1.930 ;
        RECT  2.700 1.730 3.060 1.930 ;
        RECT  2.060 0.320 3.860 0.480 ;
        RECT  3.660 0.320 3.860 1.160 ;
        RECT  3.660 0.960 4.680 1.160 ;
        RECT  2.060 0.320 2.220 1.700 ;
        RECT  1.740 1.540 2.220 1.700 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.010 2.400 ;
        RECT  3.120 1.140 6.800 2.400 ;
        RECT  0.000 1.160 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
        RECT  1.010 0.000 3.120 1.160 ;
    END
END CKMUX2M12HM

MACRO CKINVM8HM
    CLASS CORE ;
    FOREIGN CKINVM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.462  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.480 1.000 1.900 1.200 ;
        RECT  0.480 0.840 0.700 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.771  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.940 1.440 2.300 2.080 ;
        RECT  2.100 0.300 2.300 2.080 ;
        RECT  0.900 0.680 2.300 0.840 ;
        RECT  1.940 0.300 2.300 0.840 ;
        RECT  0.900 1.440 2.300 1.640 ;
        RECT  0.900 1.440 1.100 2.080 ;
        RECT  0.900 0.300 1.100 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.460 1.480 2.660 2.540 ;
        RECT  1.420 1.840 1.620 2.540 ;
        RECT  0.380 1.480 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.460 -0.140 2.660 0.580 ;
        RECT  1.380 -0.140 1.660 0.520 ;
        RECT  0.380 -0.140 0.580 0.580 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END CKINVM8HM

MACRO CKINVM6HM
    CLASS CORE ;
    FOREIGN CKINVM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.347  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.490 1.040 1.900 1.240 ;
        RECT  0.490 0.840 0.710 1.240 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.714  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 1.440 2.300 2.080 ;
        RECT  2.100 0.310 2.300 2.080 ;
        RECT  1.020 0.680 2.300 0.880 ;
        RECT  2.060 0.310 2.300 0.880 ;
        RECT  1.020 1.440 2.300 1.640 ;
        RECT  1.020 1.440 1.220 2.080 ;
        RECT  1.020 0.300 1.220 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.540 1.840 1.740 2.540 ;
        RECT  0.500 1.480 0.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.500 -0.140 1.780 0.520 ;
        RECT  0.500 -0.140 0.700 0.580 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END CKINVM6HM

MACRO CKINVM4HM
    CLASS CORE ;
    FOREIGN CKINVM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.232  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 1.100 1.280 ;
        RECT  0.100 0.840 0.300 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.386  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.740 1.440 1.500 1.640 ;
        RECT  1.300 0.680 1.500 1.640 ;
        RECT  0.740 0.680 1.500 0.840 ;
        RECT  0.740 1.440 0.940 2.080 ;
        RECT  0.740 0.300 0.940 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.260 1.840 1.460 2.540 ;
        RECT  0.220 1.480 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  1.220 -0.140 1.500 0.520 ;
        RECT  0.220 -0.140 0.420 0.580 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END CKINVM4HM

MACRO CKINVM48HM
    CLASS CORE ;
    FOREIGN CKINVM48HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 5.486  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.774  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.977  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.990 5.500 1.190 ;
        RECT  0.100 0.840 0.370 1.190 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.771  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.990 1.500 11.300 2.080 ;
        RECT  0.660 0.660 11.260 0.820 ;
        RECT  11.060 0.340 11.260 0.820 ;
        RECT  0.610 1.500 11.300 1.700 ;
        RECT  10.020 1.500 10.220 2.080 ;
        RECT  10.020 0.320 10.220 0.820 ;
        RECT  8.980 1.500 9.180 2.080 ;
        RECT  8.980 0.320 9.180 0.820 ;
        RECT  7.940 1.500 8.140 2.080 ;
        RECT  7.940 0.320 8.140 0.820 ;
        RECT  6.900 1.500 7.100 2.080 ;
        RECT  6.900 0.320 7.100 0.820 ;
        RECT  5.860 0.320 6.060 2.080 ;
        RECT  5.700 0.660 6.060 1.700 ;
        RECT  4.820 1.500 5.020 2.080 ;
        RECT  4.820 0.320 5.020 0.820 ;
        RECT  3.780 1.500 3.980 2.080 ;
        RECT  3.780 0.320 3.980 0.820 ;
        RECT  2.740 1.500 2.940 2.080 ;
        RECT  2.740 0.320 2.940 0.820 ;
        RECT  1.700 1.500 1.900 2.080 ;
        RECT  1.700 0.320 1.900 0.820 ;
        RECT  0.610 1.500 0.900 2.080 ;
        RECT  0.660 0.320 0.860 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  10.500 1.900 10.780 2.540 ;
        RECT  9.460 1.900 9.740 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  10.500 -0.140 10.780 0.500 ;
        RECT  9.460 -0.140 9.740 0.500 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  6.360 0.990 10.960 1.190 ;
        LAYER VTPH ;
        RECT  0.400 1.020 10.980 2.400 ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.020 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  10.980 0.000 11.600 1.140 ;
    END
END CKINVM48HM

MACRO CKINVM40HM
    CLASS CORE ;
    FOREIGN CKINVM40HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 4.514  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.312  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.952  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 4.700 1.200 ;
        RECT  0.100 0.840 0.310 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.863  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.940 1.500 9.220 2.080 ;
        RECT  0.660 0.680 9.180 0.840 ;
        RECT  8.980 0.320 9.180 0.840 ;
        RECT  0.620 1.500 9.220 1.700 ;
        RECT  7.940 1.500 8.140 2.080 ;
        RECT  7.940 0.320 8.140 0.840 ;
        RECT  6.900 1.500 7.100 2.080 ;
        RECT  6.900 0.320 7.100 0.840 ;
        RECT  5.860 1.500 6.060 2.080 ;
        RECT  5.860 0.320 6.060 0.840 ;
        RECT  4.900 0.680 5.200 1.700 ;
        RECT  4.820 1.500 5.020 2.080 ;
        RECT  4.820 0.320 5.020 0.840 ;
        RECT  3.780 1.500 3.980 2.080 ;
        RECT  3.780 0.320 3.980 0.840 ;
        RECT  2.740 1.500 2.940 2.080 ;
        RECT  2.740 0.320 2.940 0.840 ;
        RECT  1.700 1.500 1.900 2.080 ;
        RECT  1.700 0.320 1.900 0.840 ;
        RECT  0.620 1.500 0.900 2.080 ;
        RECT  0.660 0.320 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.500 1.480 9.700 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.500 -0.140 9.700 0.610 ;
        RECT  8.420 -0.140 8.700 0.520 ;
        RECT  7.380 -0.140 7.660 0.520 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  5.700 1.000 9.220 1.200 ;
        LAYER VTPH ;
        RECT  0.490 1.020 9.320 2.400 ;
        RECT  0.000 1.140 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.020 ;
        RECT  0.000 0.000 0.490 1.140 ;
        RECT  9.320 0.000 10.000 1.140 ;
    END
END CKINVM40HM

MACRO CKINVM3HM
    CLASS CORE ;
    FOREIGN CKINVM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.352  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.740 1.540 1.500 1.740 ;
        RECT  1.300 0.500 1.500 1.740 ;
        RECT  0.690 0.500 1.500 0.700 ;
        RECT  0.740 1.540 0.940 1.990 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 1.100 1.280 ;
        RECT  0.100 0.840 0.300 1.280 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  1.220 1.900 1.500 2.540 ;
        RECT  0.220 1.720 0.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.220 -0.140 0.420 0.670 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END CKINVM3HM

MACRO CKINVM32HM
    CLASS CORE ;
    FOREIGN CKINVM32HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 3.702  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.849  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.002  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 3.500 1.200 ;
        RECT  0.100 0.840 0.300 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.087  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.860 1.480 7.140 2.100 ;
        RECT  0.660 0.680 7.100 0.840 ;
        RECT  6.900 0.300 7.100 0.840 ;
        RECT  0.620 1.480 7.140 1.680 ;
        RECT  5.860 1.480 6.060 2.100 ;
        RECT  5.860 0.300 6.060 0.840 ;
        RECT  4.820 1.480 5.020 2.100 ;
        RECT  4.820 0.300 5.020 0.840 ;
        RECT  3.780 0.300 3.980 2.100 ;
        RECT  3.700 0.680 3.980 1.680 ;
        RECT  2.740 1.480 2.940 2.100 ;
        RECT  2.740 0.300 2.940 0.840 ;
        RECT  1.700 1.480 1.900 2.100 ;
        RECT  1.700 0.300 1.900 0.840 ;
        RECT  0.620 1.480 0.900 2.060 ;
        RECT  0.660 0.300 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.420 1.480 7.620 2.540 ;
        RECT  6.380 1.840 6.580 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        RECT  4.300 1.840 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.420 -0.140 7.620 0.610 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.160 1.000 7.320 1.200 ;
        LAYER VTPH ;
        RECT  0.450 1.020 7.310 2.400 ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.020 ;
        RECT  0.000 0.000 0.450 1.140 ;
        RECT  7.310 0.000 8.000 1.140 ;
    END
END CKINVM32HM

MACRO CKINVM2HM
    CLASS CORE ;
    FOREIGN CKINVM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.326  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.520 1.100 2.080 ;
        RECT  0.900 0.440 1.100 2.080 ;
        RECT  0.720 0.440 1.100 0.640 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.280 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.240 1.480 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.240 -0.140 0.440 0.680 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END CKINVM2HM

MACRO CKINVM24HM
    CLASS CORE ;
    FOREIGN CKINVM24HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 2.766  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.387  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.994  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 2.700 1.200 ;
        RECT  0.100 0.840 0.300 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.446  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.860 1.460 6.060 2.100 ;
        RECT  0.660 0.660 6.060 0.840 ;
        RECT  5.860 0.300 6.060 0.840 ;
        RECT  0.660 1.460 6.060 1.660 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.300 5.020 0.840 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.300 3.980 0.840 ;
        RECT  2.900 0.660 3.150 1.660 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.300 2.940 0.840 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.300 1.900 0.840 ;
        RECT  0.660 0.300 0.870 0.840 ;
        RECT  0.660 1.460 0.860 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        RECT  4.300 1.840 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.600 1.000 5.760 1.200 ;
        LAYER VTPH ;
        RECT  0.450 1.020 5.730 2.400 ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.020 ;
        RECT  0.000 0.000 0.450 1.140 ;
        RECT  5.730 0.000 6.400 1.140 ;
    END
END CKINVM24HM

MACRO CKINVM20HM
    CLASS CORE ;
    FOREIGN CKINVM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 0.998  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.156  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 0.864  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 2.300 1.220 ;
        RECT  0.100 0.840 0.300 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.069  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  0.660 0.660 5.020 0.840 ;
        RECT  4.820 0.300 5.020 0.840 ;
        RECT  0.660 1.460 5.020 1.660 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.300 3.980 0.840 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.300 2.940 0.840 ;
        RECT  2.500 0.660 2.700 1.660 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.300 1.900 0.840 ;
        RECT  0.660 1.460 0.860 2.100 ;
        RECT  0.660 0.300 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.300 1.840 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.000 1.000 4.720 1.200 ;
        LAYER VTPH ;
        RECT  0.450 1.020 4.700 2.400 ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.020 ;
        RECT  0.000 0.000 0.450 1.140 ;
        RECT  4.700 0.000 5.200 1.140 ;
    END
END CKINVM20HM

MACRO CKINVM1HM
    CLASS CORE ;
    FOREIGN CKINVM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.262  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.760 1.100 1.960 ;
        RECT  0.900 0.520 1.100 1.960 ;
        RECT  0.760 0.520 1.100 0.720 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 1.120 0.700 1.560 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.200 2.540 ;
        RECT  0.240 1.760 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.200 0.140 ;
        RECT  0.200 -0.140 0.400 0.760 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 1.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.200 1.140 ;
    END
END CKINVM1HM

MACRO CKINVM16HM
    CLASS CORE ;
    FOREIGN CKINVM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.830  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.924  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.981  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 1.900 1.200 ;
        RECT  0.100 0.840 0.360 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.540  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  0.660 0.680 3.980 0.840 ;
        RECT  3.780 0.300 3.980 0.840 ;
        RECT  0.660 1.460 3.980 1.660 ;
        RECT  2.740 1.460 2.940 2.100 ;
        RECT  2.740 0.300 2.940 0.840 ;
        RECT  2.450 0.680 2.700 1.660 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  1.700 0.300 1.900 0.840 ;
        RECT  0.660 1.460 0.860 2.100 ;
        RECT  0.660 0.300 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.300 1.480 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.300 -0.140 4.500 0.580 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.900 1.000 4.060 1.200 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END CKINVM16HM

MACRO CKINVM12HM
    CLASS CORE ;
    FOREIGN CKINVM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1.508  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.694  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.174  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 1.440 1.200 ;
        RECT  0.100 0.840 0.300 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.158  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.440 2.940 2.080 ;
        RECT  0.660 0.680 2.940 0.840 ;
        RECT  2.740 0.300 2.940 0.840 ;
        RECT  0.660 1.440 2.940 1.640 ;
        RECT  1.700 0.300 1.900 2.080 ;
        RECT  0.660 1.440 0.860 2.080 ;
        RECT  0.660 0.300 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.260 1.480 3.460 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.260 -0.140 3.460 0.580 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.160 1.000 3.160 1.200 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END CKINVM12HM

MACRO CKBUFM8HM
    CLASS CORE ;
    FOREIGN CKBUFM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.155  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 1.080 1.220 ;
        RECT  0.100 0.840 0.300 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.772  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.500 3.100 2.080 ;
        RECT  2.900 0.300 3.100 2.080 ;
        RECT  1.700 0.680 3.100 0.860 ;
        RECT  2.740 0.300 3.100 0.860 ;
        RECT  1.660 1.500 3.100 1.700 ;
        RECT  1.660 1.500 1.900 2.080 ;
        RECT  1.700 0.300 1.900 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.260 1.480 3.460 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.260 -0.140 3.460 0.580 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.340 0.860 0.860 ;
        RECT  0.660 0.680 1.500 0.860 ;
        RECT  1.300 1.020 2.700 1.220 ;
        RECT  1.300 0.680 1.500 1.740 ;
        RECT  0.660 1.540 1.500 1.740 ;
        RECT  0.660 1.540 0.860 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END CKBUFM8HM

MACRO CKBUFM6HM
    CLASS CORE ;
    FOREIGN CKBUFM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.060 0.800 1.260 ;
        RECT  0.100 1.060 0.300 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.714  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 1.460 2.700 2.100 ;
        RECT  2.500 0.300 2.700 2.100 ;
        RECT  1.420 0.680 2.700 0.840 ;
        RECT  2.460 0.300 2.700 0.840 ;
        RECT  1.420 1.460 2.700 1.660 ;
        RECT  1.420 1.460 1.620 2.100 ;
        RECT  1.420 0.300 1.620 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.940 1.840 2.140 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.520 ;
        RECT  0.860 -0.140 1.140 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 0.300 0.580 0.880 ;
        RECT  0.380 0.680 1.220 0.880 ;
        RECT  1.020 1.000 2.300 1.200 ;
        RECT  1.020 0.680 1.220 1.740 ;
        RECT  0.490 1.540 1.220 1.740 ;
        RECT  0.490 1.540 0.690 1.980 ;
        RECT  0.340 1.780 0.690 1.980 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END CKBUFM6HM

MACRO CKBUFM4HM
    CLASS CORE ;
    FOREIGN CKBUFM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.077  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.160 0.880 1.360 ;
        RECT  0.100 1.160 0.300 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.384  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.500 1.520 2.300 1.720 ;
        RECT  2.100 0.680 2.300 1.720 ;
        RECT  1.540 0.680 2.300 0.880 ;
        RECT  1.500 1.520 1.780 2.100 ;
        RECT  1.540 0.300 1.740 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  2.020 1.900 2.300 2.540 ;
        RECT  0.980 1.900 1.260 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  2.020 -0.140 2.300 0.520 ;
        RECT  0.980 -0.140 1.260 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.420 0.300 0.620 0.880 ;
        RECT  0.420 0.680 1.340 0.880 ;
        RECT  1.140 1.040 1.940 1.320 ;
        RECT  1.140 0.680 1.340 1.740 ;
        RECT  0.460 1.540 1.340 1.740 ;
        RECT  0.460 1.540 0.660 2.050 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END CKBUFM4HM

MACRO CKBUFM48HM
    CLASS CORE ;
    FOREIGN CKBUFM48HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.924  LAYER ME2  ;
        ANTENNAGATEAREA 0.924  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.992  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.100 1.500 1.300 ;
        LAYER ME2 ;
        RECT  1.300 0.940 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.980 3.680 1.340 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.725  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  14.700 1.540 14.900 2.080 ;
        RECT  4.300 0.660 14.900 0.840 ;
        RECT  14.700 0.330 14.900 0.840 ;
        RECT  4.260 1.540 14.900 1.740 ;
        RECT  13.620 1.540 13.900 2.100 ;
        RECT  13.660 0.310 13.860 0.840 ;
        RECT  12.580 1.540 12.860 2.100 ;
        RECT  12.620 0.310 12.820 0.840 ;
        RECT  11.540 1.540 11.820 2.100 ;
        RECT  11.580 0.310 11.780 0.840 ;
        RECT  10.500 1.540 10.780 2.100 ;
        RECT  10.540 0.310 10.740 0.840 ;
        RECT  9.460 1.540 9.740 2.100 ;
        RECT  9.500 0.310 9.700 0.840 ;
        RECT  9.300 0.660 9.550 1.740 ;
        RECT  8.420 1.540 8.700 2.100 ;
        RECT  8.460 0.310 8.660 0.840 ;
        RECT  7.380 1.540 7.660 2.100 ;
        RECT  7.420 0.310 7.620 0.840 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  6.380 0.310 6.580 0.840 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.310 5.540 0.840 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.310 4.500 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.200 2.540 ;
        RECT  14.140 1.900 14.420 2.540 ;
        RECT  13.100 1.900 13.380 2.540 ;
        RECT  12.060 1.900 12.340 2.540 ;
        RECT  11.020 1.900 11.300 2.540 ;
        RECT  9.980 1.900 10.260 2.540 ;
        RECT  8.940 1.900 9.220 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.200 0.140 ;
        RECT  14.140 -0.140 14.420 0.500 ;
        RECT  13.100 -0.140 13.380 0.500 ;
        RECT  12.060 -0.140 12.340 0.500 ;
        RECT  11.020 -0.140 11.300 0.500 ;
        RECT  9.980 -0.140 10.260 0.500 ;
        RECT  8.940 -0.140 9.220 0.500 ;
        RECT  7.900 -0.140 8.180 0.500 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 0.340 0.820 ;
        RECT  1.180 0.320 1.380 0.820 ;
        RECT  2.220 0.320 2.420 0.820 ;
        RECT  3.260 0.320 3.460 0.820 ;
        RECT  0.140 0.660 4.080 0.820 ;
        RECT  3.880 1.000 9.100 1.200 ;
        RECT  3.880 0.660 4.080 1.740 ;
        RECT  0.140 1.540 4.080 1.740 ;
        RECT  0.140 1.540 0.340 1.980 ;
        RECT  1.140 1.540 1.420 2.100 ;
        RECT  2.180 1.540 2.460 2.100 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  10.100 1.000 14.340 1.200 ;
        LAYER VTPH ;
        RECT  0.450 1.000 14.070 2.400 ;
        RECT  0.450 1.020 14.670 2.400 ;
        RECT  0.000 1.140 15.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.200 1.000 ;
        RECT  14.070 0.000 15.200 1.020 ;
        RECT  0.000 0.000 0.450 1.140 ;
        RECT  14.670 0.000 15.200 1.140 ;
    END
END CKBUFM48HM

MACRO CKBUFM40HM
    CLASS CORE ;
    FOREIGN CKBUFM40HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.773  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 3.020 1.200 ;
        RECT  0.100 0.840 0.300 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.889  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.100 1.460 12.300 2.100 ;
        RECT  3.780 0.660 12.300 0.820 ;
        RECT  12.100 0.300 12.300 0.820 ;
        RECT  3.780 1.460 12.300 1.660 ;
        RECT  11.060 1.460 11.260 2.100 ;
        RECT  11.060 0.300 11.260 0.820 ;
        RECT  10.020 1.460 10.220 2.100 ;
        RECT  10.020 0.300 10.220 0.820 ;
        RECT  8.980 1.460 9.180 2.100 ;
        RECT  8.980 0.300 9.180 0.820 ;
        RECT  7.940 1.460 8.140 2.100 ;
        RECT  7.940 0.300 8.140 0.820 ;
        RECT  7.700 0.660 7.950 1.660 ;
        RECT  6.900 1.460 7.100 2.100 ;
        RECT  6.900 0.300 7.100 0.820 ;
        RECT  5.860 1.460 6.060 2.100 ;
        RECT  5.860 0.300 6.060 0.820 ;
        RECT  4.820 1.460 5.020 2.100 ;
        RECT  4.820 0.300 5.020 0.820 ;
        RECT  3.780 1.460 3.980 2.100 ;
        RECT  3.780 0.300 3.980 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.620 1.840 12.820 2.540 ;
        RECT  11.580 1.840 11.780 2.540 ;
        RECT  10.540 1.840 10.740 2.540 ;
        RECT  9.500 1.840 9.700 2.540 ;
        RECT  8.460 1.840 8.660 2.540 ;
        RECT  7.420 1.840 7.620 2.540 ;
        RECT  6.380 1.840 6.580 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        RECT  4.300 1.840 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.620 -0.140 12.820 0.610 ;
        RECT  11.540 -0.140 11.820 0.500 ;
        RECT  10.500 -0.140 10.780 0.500 ;
        RECT  9.460 -0.140 9.740 0.500 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.300 0.860 0.820 ;
        RECT  1.700 0.300 1.900 0.820 ;
        RECT  2.740 0.300 2.940 0.820 ;
        RECT  0.660 0.660 3.560 0.820 ;
        RECT  3.360 0.980 7.500 1.180 ;
        RECT  3.360 0.660 3.560 1.680 ;
        RECT  0.620 1.480 3.560 1.680 ;
        RECT  0.620 1.480 0.900 2.100 ;
        RECT  1.660 1.480 1.940 2.100 ;
        RECT  2.700 1.480 2.980 2.100 ;
        RECT  8.500 0.980 12.380 1.180 ;
        LAYER VTPH ;
        RECT  0.410 1.020 12.570 2.400 ;
        RECT  0.000 1.140 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.020 ;
        RECT  0.000 0.000 0.410 1.140 ;
        RECT  12.570 0.000 13.200 1.140 ;
    END
END CKBUFM40HM

MACRO CKBUFM3HM
    CLASS CORE ;
    FOREIGN CKBUFM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.064  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.900 0.760 1.240 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.369  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.240 1.540 1.900 1.740 ;
        RECT  1.700 0.660 1.900 1.740 ;
        RECT  1.260 0.660 1.900 0.860 ;
        RECT  1.260 0.480 1.460 0.860 ;
        RECT  1.240 1.540 1.400 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.700 1.900 1.980 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  0.600 -0.140 0.880 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.540 1.080 0.740 ;
        RECT  0.920 1.060 1.500 1.260 ;
        RECT  0.920 0.540 1.080 1.740 ;
        RECT  0.180 1.540 1.080 1.740 ;
        RECT  0.180 1.540 0.380 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END CKBUFM3HM

MACRO CKBUFM32HM
    CLASS CORE ;
    FOREIGN CKBUFM32HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.614  LAYER ME1  ;
        ANTENNAGATEAREA 0.614  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.107  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.050 1.500 1.250 ;
        LAYER ME2 ;
        RECT  1.300 0.970 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.990 2.700 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.460 1.440 9.740 2.080 ;
        RECT  3.260 0.660 9.700 0.830 ;
        RECT  9.500 0.310 9.700 0.830 ;
        RECT  3.260 1.440 9.740 1.640 ;
        RECT  8.460 1.440 8.660 2.080 ;
        RECT  8.460 0.310 8.660 0.830 ;
        RECT  7.420 1.440 7.620 2.080 ;
        RECT  7.420 0.310 7.620 0.830 ;
        RECT  6.380 1.440 6.580 2.080 ;
        RECT  6.380 0.310 6.580 0.830 ;
        RECT  6.100 0.660 6.400 1.640 ;
        RECT  5.340 1.440 5.540 2.080 ;
        RECT  5.340 0.310 5.540 0.830 ;
        RECT  4.300 1.440 4.500 2.080 ;
        RECT  4.300 0.310 4.500 0.830 ;
        RECT  3.260 1.440 3.460 2.080 ;
        RECT  3.260 0.310 3.460 0.830 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.400 2.540 ;
        RECT  10.020 1.480 10.220 2.540 ;
        RECT  8.980 1.840 9.180 2.540 ;
        RECT  7.940 1.840 8.140 2.540 ;
        RECT  6.900 1.840 7.100 2.540 ;
        RECT  5.860 1.840 6.060 2.540 ;
        RECT  4.820 1.840 5.020 2.540 ;
        RECT  3.780 1.840 3.980 2.540 ;
        RECT  2.740 1.840 2.940 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.400 0.140 ;
        RECT  9.980 -0.140 10.260 0.500 ;
        RECT  8.940 -0.140 9.220 0.500 ;
        RECT  7.900 -0.140 8.180 0.500 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 0.340 0.830 ;
        RECT  1.180 0.300 1.380 0.830 ;
        RECT  2.220 0.300 2.420 0.830 ;
        RECT  0.140 0.660 3.060 0.830 ;
        RECT  2.860 0.990 5.900 1.190 ;
        RECT  2.860 0.660 3.060 1.640 ;
        RECT  0.140 1.440 3.060 1.640 ;
        RECT  0.140 1.440 0.340 2.080 ;
        RECT  1.180 1.440 1.380 2.080 ;
        RECT  2.220 1.440 2.420 2.080 ;
        RECT  6.890 0.990 9.750 1.190 ;
        LAYER VTPH ;
        RECT  1.180 1.000 9.820 2.400 ;
        RECT  0.000 1.140 10.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.400 1.000 ;
        RECT  0.000 0.000 1.180 1.140 ;
        RECT  9.820 0.000 10.400 1.140 ;
    END
END CKBUFM32HM

MACRO CKBUFM2HM
    CLASS CORE ;
    FOREIGN CKBUFM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.064  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.900 0.760 1.260 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.326  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.550 1.500 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  0.680 1.900 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.620 -0.140 0.820 0.380 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.540 1.120 0.740 ;
        RECT  0.920 0.540 1.120 1.740 ;
        RECT  0.180 1.560 1.120 1.740 ;
        RECT  0.180 1.560 0.380 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END CKBUFM2HM

MACRO CKBUFM24HM
    CLASS CORE ;
    FOREIGN CKBUFM24HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.462  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.000 2.180 1.160 ;
        RECT  0.100 0.800 0.300 1.160 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.460  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.940 1.430 8.140 2.100 ;
        RECT  2.740 0.680 8.140 0.840 ;
        RECT  7.940 0.330 8.140 0.840 ;
        RECT  2.740 1.440 8.140 1.640 ;
        RECT  5.300 1.430 8.140 1.640 ;
        RECT  6.900 1.430 7.100 2.080 ;
        RECT  6.900 0.300 7.100 0.840 ;
        RECT  5.860 1.430 6.060 2.080 ;
        RECT  5.860 0.300 6.060 0.840 ;
        RECT  5.300 0.680 5.500 1.640 ;
        RECT  4.820 1.440 5.020 2.080 ;
        RECT  4.820 0.300 5.020 0.840 ;
        RECT  3.780 1.440 3.980 2.080 ;
        RECT  3.780 0.300 3.980 0.840 ;
        RECT  2.740 1.440 2.940 2.080 ;
        RECT  2.740 0.300 2.940 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.420 1.840 7.620 2.540 ;
        RECT  6.380 1.840 6.580 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        RECT  4.300 1.840 4.500 2.540 ;
        RECT  3.260 1.840 3.460 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.380 -0.140 7.660 0.520 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.300 0.860 0.840 ;
        RECT  1.700 0.300 1.900 0.840 ;
        RECT  0.660 0.680 2.540 0.840 ;
        RECT  2.340 1.000 5.100 1.200 ;
        RECT  2.340 0.680 2.540 1.720 ;
        RECT  0.620 1.500 2.540 1.720 ;
        RECT  0.620 1.500 0.860 2.080 ;
        RECT  1.700 1.500 1.900 2.080 ;
        RECT  6.100 1.000 7.820 1.200 ;
        LAYER VTPH ;
        RECT  2.000 1.070 7.750 2.400 ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.070 ;
        RECT  0.000 0.000 2.000 1.140 ;
        RECT  7.750 0.000 8.400 1.140 ;
    END
END CKBUFM24HM

MACRO CKBUFM20HM
    CLASS CORE ;
    FOREIGN CKBUFM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.384  LAYER ME2  ;
        ANTENNAGATEAREA 0.384  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.801  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.050 1.100 1.250 ;
        LAYER ME2 ;
        RECT  0.900 0.990 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.500 0.990 1.520 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 1.440 6.620 2.080 ;
        RECT  2.220 0.660 6.580 0.840 ;
        RECT  6.380 0.310 6.580 0.840 ;
        RECT  2.220 1.440 6.620 1.640 ;
        RECT  5.340 1.440 5.540 2.080 ;
        RECT  5.340 0.300 5.540 0.840 ;
        RECT  4.300 1.440 4.500 2.080 ;
        RECT  4.300 0.300 4.500 0.840 ;
        RECT  4.100 0.660 4.350 1.640 ;
        RECT  3.260 1.440 3.460 2.080 ;
        RECT  3.260 0.300 3.460 0.840 ;
        RECT  2.220 1.440 2.420 2.080 ;
        RECT  2.220 0.310 2.420 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.860 1.840 6.060 2.540 ;
        RECT  4.820 1.840 5.020 2.540 ;
        RECT  3.780 1.840 3.980 2.540 ;
        RECT  2.740 1.840 2.940 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.310 0.340 0.830 ;
        RECT  1.180 0.300 1.380 0.830 ;
        RECT  0.140 0.660 2.000 0.830 ;
        RECT  1.820 1.000 3.900 1.200 ;
        RECT  1.820 0.660 2.000 1.660 ;
        RECT  0.140 1.460 2.000 1.660 ;
        RECT  1.180 1.460 1.380 2.080 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  4.900 1.000 6.260 1.200 ;
        LAYER VTPH ;
        RECT  0.440 1.030 6.200 2.400 ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.030 ;
        RECT  0.000 0.000 0.440 1.140 ;
        RECT  6.200 0.000 6.800 1.140 ;
    END
END CKBUFM20HM

MACRO CKBUFM1HM
    CLASS CORE ;
    FOREIGN CKBUFM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.064  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.840 0.700 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.267  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.240 0.530 1.500 2.010 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  0.700 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.620 -0.140 0.900 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.480 1.080 0.680 ;
        RECT  0.880 0.480 1.080 1.680 ;
        RECT  0.180 1.480 1.080 1.680 ;
        RECT  0.180 1.480 0.380 2.070 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END CKBUFM1HM

MACRO CKBUFM16HM
    CLASS CORE ;
    FOREIGN CKBUFM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.310  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.000 1.840 1.200 ;
        RECT  0.500 0.840 0.700 1.200 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.681  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.620 1.440 5.900 2.080 ;
        RECT  2.540 0.660 5.860 0.820 ;
        RECT  5.660 0.320 5.860 0.820 ;
        RECT  2.540 1.440 5.900 1.640 ;
        RECT  4.620 1.440 4.820 2.080 ;
        RECT  4.620 0.310 4.820 0.820 ;
        RECT  3.700 0.660 3.950 1.640 ;
        RECT  3.580 1.440 3.780 2.080 ;
        RECT  3.580 0.310 3.780 0.820 ;
        RECT  2.540 1.440 2.740 2.080 ;
        RECT  2.540 0.310 2.740 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.140 1.840 5.340 2.540 ;
        RECT  4.100 1.840 4.300 2.540 ;
        RECT  3.060 1.840 3.260 2.540 ;
        RECT  2.020 1.840 2.220 2.540 ;
        RECT  0.980 1.840 1.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.380 0.500 ;
        RECT  4.060 -0.140 4.340 0.500 ;
        RECT  3.020 -0.140 3.300 0.500 ;
        RECT  1.980 -0.140 2.260 0.500 ;
        RECT  0.980 -0.140 1.180 0.610 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.500 0.340 1.700 0.840 ;
        RECT  1.500 0.660 2.340 0.840 ;
        RECT  2.140 0.980 3.500 1.190 ;
        RECT  2.140 0.660 2.340 1.680 ;
        RECT  0.460 1.480 2.340 1.680 ;
        RECT  0.460 1.480 0.660 2.000 ;
        RECT  1.450 1.480 1.740 2.080 ;
        RECT  4.200 0.980 5.560 1.180 ;
        LAYER VTPH ;
        RECT  1.880 1.020 5.480 2.400 ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.020 ;
        RECT  0.000 0.000 1.880 1.140 ;
        RECT  5.480 0.000 6.000 1.140 ;
    END
END CKBUFM16HM

MACRO CKBUFM12HM
    CLASS CORE ;
    FOREIGN CKBUFM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.232  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 1.080 1.220 ;
        RECT  0.100 0.840 0.300 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.156  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.740 1.500 4.020 2.080 ;
        RECT  1.700 0.680 3.980 0.860 ;
        RECT  3.780 0.300 3.980 0.860 ;
        RECT  1.660 1.500 4.020 1.700 ;
        RECT  2.740 1.500 2.940 2.080 ;
        RECT  2.740 0.300 2.940 0.860 ;
        RECT  2.500 0.680 2.750 1.700 ;
        RECT  1.660 1.500 1.940 2.080 ;
        RECT  1.700 0.300 1.900 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.300 1.480 4.500 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.300 -0.140 4.500 0.580 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.520 ;
        RECT  0.140 -0.140 0.340 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.300 0.860 0.860 ;
        RECT  0.660 0.680 1.500 0.860 ;
        RECT  1.300 1.040 2.300 1.240 ;
        RECT  1.300 0.680 1.500 1.700 ;
        RECT  0.620 1.500 1.500 1.700 ;
        RECT  0.620 1.500 0.900 2.080 ;
        RECT  3.200 1.030 4.200 1.250 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END CKBUFM12HM

MACRO CKAN2M8HM
    CLASS CORE ;
    FOREIGN CKAN2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.700 1.180 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.144  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.180 1.200 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.866  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.450 3.100 2.090 ;
        RECT  2.900 0.340 3.100 2.090 ;
        RECT  1.780 0.660 3.100 0.860 ;
        RECT  2.840 0.340 3.100 0.860 ;
        RECT  1.700 1.450 3.100 1.690 ;
        RECT  1.780 0.340 1.980 0.860 ;
        RECT  1.700 1.450 1.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.280 1.480 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.260 -0.140 2.540 0.500 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.340 0.370 0.540 0.660 ;
        RECT  0.340 0.480 1.540 0.660 ;
        RECT  1.340 1.040 2.740 1.240 ;
        RECT  1.340 0.480 1.540 1.710 ;
        RECT  0.620 1.510 1.540 1.710 ;
        RECT  0.620 1.510 0.840 2.090 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END CKAN2M8HM

MACRO CKAN2M6HM
    CLASS CORE ;
    FOREIGN CKAN2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.680 1.170 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.140  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.180 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.702  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 1.480 3.100 2.080 ;
        RECT  2.870 0.740 3.100 2.080 ;
        RECT  1.780 0.740 3.100 0.920 ;
        RECT  1.740 1.480 3.100 1.700 ;
        RECT  1.740 1.480 2.020 2.080 ;
        RECT  1.780 0.380 1.980 0.920 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.260 -0.140 2.540 0.520 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.260 0.500 1.550 0.660 ;
        RECT  1.350 1.090 2.690 1.290 ;
        RECT  1.350 0.500 1.550 1.720 ;
        RECT  0.620 1.510 1.550 1.720 ;
        RECT  0.620 1.510 0.900 2.090 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END CKAN2M6HM

MACRO CKAN2M4HM
    CLASS CORE ;
    FOREIGN CKAN2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.700 1.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.094  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.180 1.200 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.740 1.460 2.300 1.700 ;
        RECT  2.100 0.670 2.300 1.700 ;
        RECT  1.780 0.670 2.300 0.850 ;
        RECT  1.740 1.460 2.020 2.080 ;
        RECT  1.780 0.310 1.980 0.850 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.140 1.540 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.260 -0.140 2.540 0.500 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.340 0.320 0.540 0.670 ;
        RECT  0.340 0.490 1.550 0.670 ;
        RECT  1.350 1.040 1.940 1.240 ;
        RECT  1.350 0.490 1.550 1.740 ;
        RECT  0.580 1.540 1.550 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END CKAN2M4HM

MACRO CKAN2M3HM
    CLASS CORE ;
    FOREIGN CKAN2M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.170 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.067  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.830 1.100 1.190 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.413  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.600 1.430 2.300 1.720 ;
        RECT  2.100 0.360 2.300 1.720 ;
        RECT  1.680 0.360 2.300 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  2.020 2.020 2.300 2.540 ;
        RECT  0.510 2.020 0.870 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.040 -0.140 1.320 0.340 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.440 0.380 0.660 ;
        RECT  0.100 0.500 1.460 0.660 ;
        RECT  1.270 0.500 1.460 1.170 ;
        RECT  1.270 0.890 1.940 1.170 ;
        RECT  1.270 0.500 1.440 1.680 ;
        RECT  0.500 1.520 1.440 1.680 ;
        LAYER VTPH ;
        RECT  0.850 1.070 2.400 2.400 ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.070 ;
        RECT  0.000 0.000 0.850 1.140 ;
    END
END CKAN2M3HM

MACRO CKAN2M2HM
    CLASS CORE ;
    FOREIGN CKAN2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.049  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.049  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 0.840 1.140 1.200 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.340  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.460 1.900 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.100 2.000 1.300 2.540 ;
        RECT  0.140 2.000 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.040 -0.140 1.320 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.450 0.380 0.670 ;
        RECT  0.100 0.480 1.520 0.670 ;
        RECT  1.320 0.480 1.520 1.720 ;
        RECT  0.580 1.500 1.520 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END CKAN2M2HM

MACRO CKAN2M16HM
    CLASS CORE ;
    FOREIGN CKAN2M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.293  LAYER ME1  ;
        ANTENNAGATEAREA 0.293  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.669  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.160 1.500 1.360 ;
        LAYER ME2 ;
        RECT  1.300 1.020 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.910 1.120 1.570 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.293  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.860 0.800 2.060 1.180 ;
        RECT  0.440 0.800 2.060 0.960 ;
        RECT  0.440 0.800 0.700 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.684  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.880 1.500 6.100 2.080 ;
        RECT  2.700 1.500 6.100 1.700 ;
        RECT  4.820 1.500 5.020 2.080 ;
        RECT  2.740 0.660 5.020 0.860 ;
        RECT  4.820 0.370 5.020 0.860 ;
        RECT  4.100 0.660 4.350 1.700 ;
        RECT  3.780 1.500 3.980 2.080 ;
        RECT  3.780 0.370 3.980 0.860 ;
        RECT  2.700 1.500 2.960 2.080 ;
        RECT  2.740 0.380 2.940 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.380 1.470 6.580 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.080 -0.140 2.360 0.320 ;
        RECT  0.260 -0.140 0.460 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.080 0.480 2.440 0.640 ;
        RECT  2.240 1.070 3.940 1.270 ;
        RECT  2.240 0.480 2.440 1.740 ;
        RECT  0.620 1.580 2.440 1.740 ;
        RECT  1.700 1.580 1.900 2.050 ;
        RECT  0.620 1.580 0.840 2.060 ;
        RECT  4.860 1.070 6.220 1.270 ;
        LAYER VTPH ;
        RECT  0.750 1.100 2.600 2.400 ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.100 ;
        RECT  0.000 0.000 0.750 1.140 ;
        RECT  2.600 0.000 6.800 1.140 ;
    END
END CKAN2M16HM

MACRO CKAN2M12HM
    CLASS CORE ;
    FOREIGN CKAN2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.282  LAYER ME1  ;
        ANTENNAGATEAREA 0.282  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.678  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 1.000 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.950 1.120 1.620 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.282  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.820 0.800 2.100 1.150 ;
        RECT  0.100 0.800 2.100 0.960 ;
        RECT  0.100 0.800 0.760 1.160 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.208  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.840 1.500 5.060 2.080 ;
        RECT  2.700 1.500 5.060 1.700 ;
        RECT  3.780 0.380 3.980 2.080 ;
        RECT  3.700 0.680 3.980 1.700 ;
        RECT  2.740 0.680 3.980 0.880 ;
        RECT  2.740 0.380 2.940 0.880 ;
        RECT  2.700 1.500 2.920 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.340 1.460 5.540 2.540 ;
        RECT  4.260 1.880 4.540 2.540 ;
        RECT  3.220 1.880 3.500 2.540 ;
        RECT  2.180 1.880 2.460 2.540 ;
        RECT  1.140 1.880 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.080 -0.140 2.360 0.320 ;
        RECT  0.100 -0.140 0.380 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.100 0.480 2.500 0.640 ;
        RECT  2.300 1.080 3.540 1.280 ;
        RECT  2.300 0.480 2.500 1.700 ;
        RECT  0.620 1.540 2.500 1.700 ;
        RECT  0.620 1.540 0.890 2.020 ;
        RECT  1.660 1.540 1.940 2.020 ;
        RECT  4.460 1.080 5.260 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END CKAN2M12HM

MACRO BUFTM8HM
    CLASS CORE ;
    FOREIGN BUFTM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.173  LAYER ME1  ;
        ANTENNAGATEAREA 0.173  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 0.990 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.080 0.700 1.400 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.050 2.770 1.560 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.069  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.120 0.900 5.860 1.100 ;
        RECT  5.660 0.340 5.860 1.100 ;
        RECT  5.140 0.900 5.340 2.100 ;
        RECT  4.120 0.680 4.770 1.100 ;
        RECT  4.570 0.350 4.770 1.100 ;
        RECT  4.120 0.680 4.300 2.030 ;
        RECT  3.530 0.680 4.770 0.880 ;
        RECT  3.530 0.350 3.730 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.660 1.480 5.860 2.540 ;
        RECT  4.620 1.480 4.820 2.540 ;
        RECT  3.510 1.870 3.790 2.540 ;
        RECT  2.400 2.080 2.680 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.090 -0.140 5.290 0.580 ;
        RECT  4.010 -0.140 4.290 0.520 ;
        RECT  2.930 -0.140 3.210 0.320 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.310 0.320 0.860 ;
        RECT  0.160 0.700 1.040 0.860 ;
        RECT  0.880 0.700 1.040 1.720 ;
        RECT  0.160 1.560 1.040 1.720 ;
        RECT  0.160 1.560 0.320 2.100 ;
        RECT  1.240 0.300 2.610 0.460 ;
        RECT  2.410 0.300 2.610 0.700 ;
        RECT  2.410 0.500 3.370 0.700 ;
        RECT  3.170 0.500 3.370 1.110 ;
        RECT  1.240 0.300 1.400 1.590 ;
        RECT  1.240 1.430 1.920 1.590 ;
        RECT  1.700 1.430 1.920 1.770 ;
        RECT  1.740 0.620 2.240 0.780 ;
        RECT  3.760 1.160 3.960 1.710 ;
        RECT  2.960 1.550 3.960 1.710 ;
        RECT  2.960 1.550 3.240 1.920 ;
        RECT  2.080 1.730 3.240 1.920 ;
        RECT  1.180 1.820 1.380 2.100 ;
        RECT  2.080 0.620 2.240 2.100 ;
        RECT  1.180 1.940 2.240 2.100 ;
        LAYER VTPH ;
        RECT  3.330 1.070 5.480 2.400 ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.580 1.190 2.250 2.400 ;
        RECT  0.000 1.210 2.250 2.400 ;
        RECT  3.330 1.140 6.000 2.400 ;
        RECT  0.000 1.320 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.070 ;
        RECT  0.000 0.000 3.330 1.140 ;
        RECT  5.480 0.000 6.000 1.140 ;
        RECT  0.400 0.000 3.330 1.190 ;
        RECT  0.400 0.000 1.580 1.210 ;
        RECT  2.250 0.000 3.330 1.320 ;
    END
END BUFTM8HM

MACRO BUFTM6HM
    CLASS CORE ;
    FOREIGN BUFTM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.761  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.060 2.700 1.260 ;
        LAYER ME2 ;
        RECT  2.500 0.990 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.470 1.000 2.870 1.390 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.166  LAYER ME1  ;
        ANTENNAGATEAREA 0.166  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 0.990 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.080 0.700 1.400 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.744  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.490 1.570 4.700 2.030 ;
        RECT  4.500 0.310 4.700 2.030 ;
        RECT  3.470 0.680 4.700 0.880 ;
        RECT  4.490 0.310 4.700 0.880 ;
        RECT  3.450 1.570 4.700 1.740 ;
        RECT  3.450 1.570 3.650 2.030 ;
        RECT  3.470 0.310 3.630 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.010 1.710 5.210 2.540 ;
        RECT  3.930 1.900 4.210 2.540 ;
        RECT  2.860 1.870 3.140 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.010 -0.140 5.210 0.630 ;
        RECT  3.930 -0.140 4.210 0.520 ;
        RECT  2.860 -0.140 3.140 0.520 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.350 0.340 0.860 ;
        RECT  0.140 0.700 1.040 0.860 ;
        RECT  0.880 0.700 1.040 1.720 ;
        RECT  0.140 1.560 1.040 1.720 ;
        RECT  0.140 1.560 0.340 2.060 ;
        RECT  1.240 0.300 2.530 0.460 ;
        RECT  2.370 0.300 2.530 0.840 ;
        RECT  2.370 0.680 3.310 0.840 ;
        RECT  3.110 0.680 3.310 1.080 ;
        RECT  1.240 0.300 1.400 1.590 ;
        RECT  1.240 1.430 1.980 1.590 ;
        RECT  1.700 1.430 1.980 1.780 ;
        RECT  1.740 0.620 2.100 0.780 ;
        RECT  1.940 0.620 2.100 1.240 ;
        RECT  1.940 1.080 2.310 1.240 ;
        RECT  3.130 1.250 3.870 1.410 ;
        RECT  2.150 1.080 2.310 1.710 ;
        RECT  3.130 1.250 3.290 1.710 ;
        RECT  2.150 1.550 3.290 1.710 ;
        RECT  1.180 1.820 1.380 2.100 ;
        RECT  2.370 1.550 2.530 2.100 ;
        RECT  1.180 1.940 2.530 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.800 1.140 5.600 2.400 ;
        RECT  0.000 1.210 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
        RECT  0.400 0.000 1.800 1.210 ;
    END
END BUFTM6HM

MACRO BUFTM4HM
    CLASS CORE ;
    FOREIGN BUFTM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.663  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.120 2.700 1.320 ;
        LAYER ME2 ;
        RECT  2.500 1.010 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.000 2.780 1.390 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.166  LAYER ME1  ;
        ANTENNAGATEAREA 0.166  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.575  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 1.010 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.080 0.700 1.400 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.608  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.380 0.330 4.580 2.030 ;
        RECT  3.340 1.300 4.580 1.500 ;
        RECT  3.340 0.330 3.540 2.020 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.860 1.750 4.060 2.540 ;
        RECT  2.780 1.870 3.060 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.860 -0.140 4.060 0.600 ;
        RECT  2.780 -0.140 3.060 0.520 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.310 0.320 0.860 ;
        RECT  0.160 0.700 1.040 0.860 ;
        RECT  0.880 0.700 1.040 1.720 ;
        RECT  0.160 1.560 1.040 1.720 ;
        RECT  0.160 1.560 0.320 2.100 ;
        RECT  1.740 0.620 2.100 0.780 ;
        RECT  1.940 0.620 2.100 1.240 ;
        RECT  1.940 1.080 2.300 1.240 ;
        RECT  2.140 1.080 2.300 1.710 ;
        RECT  2.940 1.280 3.140 1.710 ;
        RECT  2.140 1.550 3.140 1.710 ;
        RECT  1.200 1.750 1.420 2.100 ;
        RECT  2.320 1.550 2.480 2.100 ;
        RECT  1.200 1.940 2.480 2.100 ;
        RECT  1.240 0.300 2.500 0.460 ;
        RECT  2.300 0.300 2.500 0.840 ;
        RECT  2.300 0.680 3.160 0.840 ;
        RECT  2.960 0.680 3.160 1.040 ;
        RECT  1.240 0.300 1.400 1.590 ;
        RECT  1.240 1.430 1.980 1.590 ;
        RECT  1.700 1.430 1.980 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.800 1.140 4.800 2.400 ;
        RECT  0.000 1.210 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
        RECT  0.400 0.000 1.800 1.210 ;
    END
END BUFTM4HM

MACRO BUFTM3HM
    CLASS CORE ;
    FOREIGN BUFTM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.459  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.700 1.120 2.900 1.320 ;
        LAYER ME1 ;
        RECT  2.660 1.000 2.980 1.390 ;
        LAYER ME2 ;
        RECT  2.700 1.010 3.100 1.560 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.166  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.090 0.760 1.290 ;
        RECT  0.100 0.800 0.300 1.290 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.412  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.540 1.150 3.900 1.560 ;
        RECT  3.540 0.330 3.740 2.020 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  4.060 1.750 4.260 2.540 ;
        RECT  2.980 1.870 3.260 2.540 ;
        RECT  0.820 1.900 1.100 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  4.060 -0.140 4.260 0.600 ;
        RECT  2.980 -0.140 3.260 0.520 ;
        RECT  0.820 -0.140 1.100 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.300 0.360 0.640 0.560 ;
        RECT  0.480 0.360 0.640 0.860 ;
        RECT  0.480 0.700 1.240 0.860 ;
        RECT  1.080 0.700 1.240 1.720 ;
        RECT  0.360 1.560 1.240 1.720 ;
        RECT  0.360 1.560 0.520 2.100 ;
        RECT  1.980 0.620 2.270 1.240 ;
        RECT  1.980 1.040 2.500 1.240 ;
        RECT  2.340 1.040 2.500 1.710 ;
        RECT  3.140 1.240 3.340 1.710 ;
        RECT  2.340 1.550 3.340 1.710 ;
        RECT  1.400 1.750 1.620 2.100 ;
        RECT  2.520 1.550 2.680 2.100 ;
        RECT  1.400 1.940 2.680 2.100 ;
        RECT  1.440 0.300 2.740 0.460 ;
        RECT  2.470 0.300 2.740 0.840 ;
        RECT  2.470 0.680 3.340 0.840 ;
        RECT  3.140 0.680 3.340 1.010 ;
        RECT  1.440 0.300 1.600 1.590 ;
        RECT  1.440 1.430 2.180 1.590 ;
        RECT  1.900 1.430 2.180 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.600 2.400 ;
        RECT  2.000 1.140 4.400 2.400 ;
        RECT  0.000 1.210 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
        RECT  0.600 0.000 2.000 1.210 ;
    END
END BUFTM3HM

MACRO BUFTM2HM
    CLASS CORE ;
    FOREIGN BUFTM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.166  LAYER ME1  ;
        ANTENNAGATEAREA 0.166  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 1.010 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.080 0.700 1.400 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.145  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.120 2.700 1.320 ;
        LAYER ME2 ;
        RECT  2.500 1.010 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.050 2.780 1.390 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.270 1.440 3.900 2.080 ;
        RECT  3.740 0.310 3.900 2.080 ;
        RECT  3.580 0.310 3.900 0.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  2.700 1.870 2.980 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.940 -0.140 3.220 0.500 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.320 0.340 0.860 ;
        RECT  0.140 0.700 1.040 0.860 ;
        RECT  0.880 0.700 1.040 1.720 ;
        RECT  0.160 1.560 1.040 1.720 ;
        RECT  0.160 1.560 0.320 2.100 ;
        RECT  1.780 0.620 2.070 1.240 ;
        RECT  1.780 1.040 2.300 1.240 ;
        RECT  2.140 1.040 2.300 2.100 ;
        RECT  2.940 1.020 3.100 1.710 ;
        RECT  2.140 1.550 3.100 1.710 ;
        RECT  1.180 1.820 1.380 2.100 ;
        RECT  2.140 1.550 2.400 2.100 ;
        RECT  1.180 1.940 2.400 2.100 ;
        RECT  1.240 0.300 2.560 0.460 ;
        RECT  2.360 0.300 2.560 0.850 ;
        RECT  2.360 0.690 3.580 0.850 ;
        RECT  3.360 0.690 3.580 1.220 ;
        RECT  1.240 0.300 1.400 1.590 ;
        RECT  1.240 1.430 1.980 1.590 ;
        RECT  1.700 1.430 1.980 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.800 1.140 4.000 2.400 ;
        RECT  0.000 1.210 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  0.400 0.000 1.800 1.210 ;
    END
END BUFTM2HM

MACRO BUFTM24HM
    CLASS CORE ;
    FOREIGN BUFTM24HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.599  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.040 4.700 1.240 ;
        LAYER ME2 ;
        RECT  4.500 0.840 4.700 1.560 ;
        LAYER ME1 ;
        RECT  3.520 1.010 5.080 1.280 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.324  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.790 0.360 1.360 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.864  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.410 1.490 11.700 2.100 ;
        RECT  6.300 0.660 11.700 0.820 ;
        RECT  11.500 0.390 11.700 0.820 ;
        RECT  6.260 1.510 11.700 1.720 ;
        RECT  8.800 1.490 11.700 1.720 ;
        RECT  10.380 1.490 10.660 2.080 ;
        RECT  10.460 0.390 10.660 0.820 ;
        RECT  9.330 1.490 9.630 2.090 ;
        RECT  9.420 0.390 9.620 0.820 ;
        RECT  8.800 0.660 9.150 1.720 ;
        RECT  8.300 1.510 8.580 2.090 ;
        RECT  8.380 0.390 8.580 0.820 ;
        RECT  7.250 1.510 7.560 2.090 ;
        RECT  7.340 0.390 7.540 0.820 ;
        RECT  6.260 1.510 7.560 1.740 ;
        RECT  6.300 0.390 6.500 0.820 ;
        RECT  6.260 1.510 6.460 2.030 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.400 2.540 ;
        RECT  11.980 1.480 12.180 2.540 ;
        RECT  10.900 1.900 11.180 2.540 ;
        RECT  9.860 1.900 10.140 2.540 ;
        RECT  8.820 1.900 9.100 2.540 ;
        RECT  7.780 1.900 8.060 2.540 ;
        RECT  6.740 1.900 7.020 2.540 ;
        RECT  5.660 1.950 5.940 2.540 ;
        RECT  4.780 1.880 5.060 2.540 ;
        RECT  3.740 1.880 4.020 2.540 ;
        RECT  1.740 2.020 1.980 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.400 0.140 ;
        RECT  12.020 -0.140 12.220 0.630 ;
        RECT  10.940 -0.140 11.220 0.500 ;
        RECT  9.900 -0.140 10.180 0.500 ;
        RECT  8.860 -0.140 9.140 0.500 ;
        RECT  7.820 -0.140 8.100 0.500 ;
        RECT  6.780 -0.140 7.060 0.500 ;
        RECT  5.740 -0.140 6.020 0.500 ;
        RECT  4.740 -0.140 5.020 0.500 ;
        RECT  3.700 -0.140 3.980 0.500 ;
        RECT  2.660 -0.140 2.940 0.500 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.300 0.860 0.870 ;
        RECT  0.660 0.660 1.200 0.870 ;
        RECT  1.020 1.330 2.150 1.500 ;
        RECT  1.020 0.660 1.200 1.720 ;
        RECT  0.140 1.560 1.200 1.720 ;
        RECT  0.140 1.560 0.340 2.080 ;
        RECT  1.100 0.300 2.360 0.460 ;
        RECT  1.100 0.300 1.400 0.500 ;
        RECT  2.200 0.300 2.360 0.820 ;
        RECT  3.220 0.310 3.420 0.840 ;
        RECT  4.260 0.390 4.460 0.840 ;
        RECT  2.200 0.660 5.540 0.820 ;
        RECT  5.250 0.310 5.540 0.840 ;
        RECT  2.760 0.700 5.780 0.840 ;
        RECT  5.280 0.700 5.780 0.900 ;
        RECT  2.760 0.660 2.960 1.780 ;
        RECT  1.610 0.620 1.910 1.160 ;
        RECT  1.610 0.990 2.600 1.160 ;
        RECT  5.800 1.200 6.080 1.720 ;
        RECT  3.220 1.480 6.080 1.720 ;
        RECT  1.380 1.680 2.600 1.860 ;
        RECT  2.440 0.990 2.600 2.100 ;
        RECT  1.380 1.680 1.560 2.080 ;
        RECT  1.140 1.880 1.560 2.080 ;
        RECT  4.260 1.480 4.530 2.090 ;
        RECT  3.220 1.480 3.500 2.100 ;
        RECT  2.440 1.940 3.500 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 12.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.400 1.140 ;
    END
END BUFTM24HM

MACRO BUFTM20HM
    CLASS CORE ;
    FOREIGN BUFTM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.500  LAYER ME1  ;
        ANTENNAGATEAREA 0.500  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.756  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.160 4.700 1.360 ;
        LAYER ME2 ;
        RECT  4.500 1.010 4.700 1.560 ;
        LAYER ME1 ;
        RECT  3.530 1.120 4.960 1.380 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.287  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.790 0.420 1.250 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.500  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.700 1.450 10.980 2.080 ;
        RECT  6.580 0.660 10.940 0.890 ;
        RECT  10.740 0.390 10.940 0.890 ;
        RECT  6.590 1.470 10.980 1.720 ;
        RECT  9.250 1.450 10.980 1.720 ;
        RECT  9.650 1.450 9.950 2.090 ;
        RECT  9.700 0.390 9.900 0.890 ;
        RECT  9.250 0.660 9.550 1.720 ;
        RECT  8.620 1.470 8.900 2.090 ;
        RECT  8.660 0.390 8.860 0.890 ;
        RECT  7.570 1.470 7.880 2.090 ;
        RECT  7.620 0.390 7.820 0.890 ;
        RECT  6.590 1.470 7.880 1.740 ;
        RECT  6.590 1.470 6.780 2.050 ;
        RECT  6.580 0.390 6.780 0.890 ;
        RECT  5.470 0.480 6.780 0.640 ;
        RECT  5.470 0.330 5.690 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.260 1.480 11.460 2.540 ;
        RECT  10.180 1.900 10.460 2.540 ;
        RECT  9.140 1.900 9.420 2.540 ;
        RECT  8.100 1.900 8.380 2.540 ;
        RECT  7.060 1.900 7.340 2.540 ;
        RECT  6.020 1.900 6.320 2.540 ;
        RECT  4.780 1.880 5.060 2.540 ;
        RECT  3.740 1.880 4.020 2.540 ;
        RECT  1.740 2.020 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.260 -0.140 11.460 0.630 ;
        RECT  10.180 -0.140 10.460 0.500 ;
        RECT  9.140 -0.140 9.420 0.500 ;
        RECT  8.100 -0.140 8.380 0.500 ;
        RECT  7.060 -0.140 7.340 0.500 ;
        RECT  5.980 -0.140 6.260 0.320 ;
        RECT  4.840 -0.140 5.120 0.500 ;
        RECT  3.790 -0.140 4.070 0.500 ;
        RECT  2.750 -0.140 3.030 0.500 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.330 2.120 1.500 ;
        RECT  0.660 0.300 0.860 1.730 ;
        RECT  0.140 1.560 0.860 1.730 ;
        RECT  0.140 1.560 0.340 2.080 ;
        RECT  1.130 0.300 2.450 0.460 ;
        RECT  2.150 0.300 2.450 0.820 ;
        RECT  3.310 0.310 3.510 0.840 ;
        RECT  4.350 0.390 4.550 0.840 ;
        RECT  1.130 0.300 1.350 0.760 ;
        RECT  2.150 0.660 5.300 0.820 ;
        RECT  2.720 0.660 5.300 0.840 ;
        RECT  5.130 0.660 5.300 1.080 ;
        RECT  5.130 0.920 5.660 1.080 ;
        RECT  2.720 0.660 2.920 1.780 ;
        RECT  1.610 0.620 1.910 1.160 ;
        RECT  1.610 0.990 2.540 1.160 ;
        RECT  5.840 1.200 6.420 1.720 ;
        RECT  3.260 1.560 6.420 1.720 ;
        RECT  1.180 1.670 2.540 1.860 ;
        RECT  2.330 0.990 2.540 2.100 ;
        RECT  2.310 1.670 2.540 2.100 ;
        RECT  4.300 1.560 4.500 2.010 ;
        RECT  5.340 1.560 5.540 2.010 ;
        RECT  1.180 1.670 1.380 2.060 ;
        RECT  3.260 1.560 3.460 2.100 ;
        RECT  2.310 1.940 3.460 2.100 ;
        LAYER VTPH ;
        RECT  5.980 1.060 11.170 2.400 ;
        RECT  0.000 1.140 3.650 2.400 ;
        RECT  5.980 1.140 11.600 2.400 ;
        RECT  0.000 1.240 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.060 ;
        RECT  0.000 0.000 5.980 1.140 ;
        RECT  11.170 0.000 11.600 1.140 ;
        RECT  3.650 0.000 5.980 1.240 ;
    END
END BUFTM20HM

MACRO BUFTM1HM
    CLASS CORE ;
    FOREIGN BUFTM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.145  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.120 2.700 1.320 ;
        LAYER ME2 ;
        RECT  2.500 1.010 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.460 1.050 2.780 1.390 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.166  LAYER ME1  ;
        ANTENNAGATEAREA 0.166  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.889  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 1.010 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.080 0.700 1.400 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 1.640 3.630 2.030 ;
        RECT  3.420 0.310 3.630 2.030 ;
        RECT  3.280 0.310 3.630 0.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  2.700 1.870 2.980 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.780 -0.140 3.060 0.500 ;
        RECT  0.620 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.320 0.340 0.860 ;
        RECT  0.140 0.700 1.040 0.860 ;
        RECT  0.880 0.700 1.040 1.720 ;
        RECT  0.160 1.560 1.040 1.720 ;
        RECT  0.160 1.560 0.320 2.100 ;
        RECT  1.780 0.620 2.060 1.240 ;
        RECT  1.780 1.040 2.300 1.240 ;
        RECT  2.140 1.040 2.300 2.100 ;
        RECT  2.940 1.220 3.100 1.710 ;
        RECT  2.140 1.550 3.100 1.710 ;
        RECT  1.200 1.750 1.420 2.100 ;
        RECT  2.140 1.550 2.400 2.100 ;
        RECT  1.200 1.940 2.400 2.100 ;
        RECT  1.240 0.300 2.500 0.460 ;
        RECT  2.300 0.300 2.500 0.850 ;
        RECT  2.300 0.690 3.200 0.850 ;
        RECT  3.000 0.690 3.200 1.050 ;
        RECT  1.240 0.300 1.400 1.590 ;
        RECT  1.240 1.430 1.980 1.590 ;
        RECT  1.700 1.430 1.980 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  1.800 1.140 4.000 2.400 ;
        RECT  0.000 1.210 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
        RECT  0.400 0.000 1.800 1.210 ;
    END
END BUFTM1HM

MACRO BUFTM16HM
    CLASS CORE ;
    FOREIGN BUFTM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.365  LAYER ME1  ;
        ANTENNAGATEAREA 0.365  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.311  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.140 3.100 1.340 ;
        LAYER ME2 ;
        RECT  2.900 1.000 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.900 1.080 3.500 1.400 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.076  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 1.000 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.080 0.700 1.400 ;
        END
    END E
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.050  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.220 0.680 8.460 0.880 ;
        RECT  8.260 0.390 8.460 0.880 ;
        RECT  7.740 1.430 7.940 2.090 ;
        RECT  5.620 1.430 7.940 1.720 ;
        RECT  7.220 0.390 7.420 0.880 ;
        RECT  6.660 1.430 6.940 2.080 ;
        RECT  6.180 0.390 6.380 0.880 ;
        RECT  6.050 0.680 6.300 1.720 ;
        RECT  5.620 1.430 5.900 2.080 ;
        RECT  4.620 1.580 5.900 1.740 ;
        RECT  5.140 0.390 5.340 0.880 ;
        RECT  4.620 1.580 4.820 1.990 ;
        RECT  4.220 0.320 4.420 0.880 ;
        RECT  4.060 0.320 4.420 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.260 1.480 8.460 2.540 ;
        RECT  7.180 1.900 7.460 2.540 ;
        RECT  6.140 1.900 6.420 2.540 ;
        RECT  5.100 1.900 5.380 2.540 ;
        RECT  4.060 1.900 4.340 2.540 ;
        RECT  3.020 1.900 3.300 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  7.700 -0.140 7.980 0.520 ;
        RECT  6.660 -0.140 6.940 0.520 ;
        RECT  5.620 -0.140 5.900 0.520 ;
        RECT  4.580 -0.140 4.860 0.520 ;
        RECT  3.540 -0.140 3.820 0.520 ;
        RECT  2.460 -0.140 2.740 0.320 ;
        RECT  0.660 -0.140 0.860 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.360 0.380 0.900 ;
        RECT  0.100 0.740 1.020 0.900 ;
        RECT  0.860 0.740 1.020 1.740 ;
        RECT  0.860 1.440 1.820 1.740 ;
        RECT  0.140 1.580 1.820 1.740 ;
        RECT  0.140 1.580 0.340 2.060 ;
        RECT  1.200 0.300 2.300 0.460 ;
        RECT  2.140 0.300 2.300 0.640 ;
        RECT  2.140 0.480 3.260 0.640 ;
        RECT  3.060 0.480 3.260 0.840 ;
        RECT  3.060 0.680 4.060 0.840 ;
        RECT  1.200 0.300 1.360 1.280 ;
        RECT  3.860 0.680 4.060 1.140 ;
        RECT  1.200 1.120 2.260 1.280 ;
        RECT  1.980 1.120 2.260 1.780 ;
        RECT  1.650 0.630 1.940 0.960 ;
        RECT  1.650 0.800 2.720 0.960 ;
        RECT  4.270 1.200 4.630 1.420 ;
        RECT  4.270 1.200 4.460 1.740 ;
        RECT  2.560 1.580 4.460 1.740 ;
        RECT  1.230 1.900 1.610 2.100 ;
        RECT  3.540 1.580 3.820 2.010 ;
        RECT  2.560 0.800 2.720 2.100 ;
        RECT  1.230 1.940 2.720 2.100 ;
        LAYER VTPH ;
        RECT  4.580 1.120 7.980 2.400 ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  3.990 1.140 8.800 2.400 ;
        RECT  0.000 1.260 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.120 ;
        RECT  0.000 0.000 4.580 1.140 ;
        RECT  7.980 0.000 8.800 1.140 ;
        RECT  0.400 0.000 3.990 1.260 ;
    END
END BUFTM16HM

MACRO BUFTM12HM
    CLASS CORE ;
    FOREIGN BUFTM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.197  LAYER ME1  ;
        ANTENNAGATEAREA 0.197  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.431  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.140 0.700 1.340 ;
        LAYER ME2 ;
        RECT  0.500 0.990 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.100 1.080 0.700 1.400 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.790 1.170 3.330 1.500 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.569  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.680 0.900 7.460 1.100 ;
        RECT  7.260 0.400 7.460 1.100 ;
        RECT  6.690 0.900 6.980 1.990 ;
        RECT  6.220 0.340 6.420 1.100 ;
        RECT  5.700 0.900 5.900 2.100 ;
        RECT  4.680 0.680 5.330 1.100 ;
        RECT  5.130 0.350 5.330 1.100 ;
        RECT  4.680 0.680 4.860 2.030 ;
        RECT  4.090 0.680 5.330 0.880 ;
        RECT  4.090 0.350 4.290 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  7.260 1.480 7.460 2.540 ;
        RECT  6.220 1.480 6.420 2.540 ;
        RECT  5.180 1.480 5.380 2.540 ;
        RECT  4.070 1.870 4.350 2.540 ;
        RECT  2.960 2.080 3.240 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.740 -0.140 6.940 0.580 ;
        RECT  5.650 -0.140 5.850 0.580 ;
        RECT  4.570 -0.140 4.850 0.520 ;
        RECT  3.570 -0.140 3.770 0.560 ;
        RECT  2.490 -0.140 2.690 0.560 ;
        RECT  0.600 -0.140 0.900 0.540 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.310 0.320 0.860 ;
        RECT  0.160 0.700 1.040 0.860 ;
        RECT  0.880 0.700 1.040 1.720 ;
        RECT  0.160 1.560 1.040 1.720 ;
        RECT  0.160 1.560 0.320 2.100 ;
        RECT  1.240 0.300 2.320 0.460 ;
        RECT  2.160 0.300 2.320 0.910 ;
        RECT  3.010 0.440 3.210 0.910 ;
        RECT  2.160 0.750 3.930 0.910 ;
        RECT  3.730 0.750 3.930 1.150 ;
        RECT  1.240 0.300 1.400 1.590 ;
        RECT  1.240 1.430 1.980 1.590 ;
        RECT  1.700 1.430 1.980 1.780 ;
        RECT  1.780 0.640 2.000 1.230 ;
        RECT  1.780 1.070 2.300 1.230 ;
        RECT  4.280 1.180 4.500 1.710 ;
        RECT  3.520 1.550 4.500 1.710 ;
        RECT  3.520 1.550 3.800 1.920 ;
        RECT  2.140 1.760 3.800 1.920 ;
        RECT  1.180 1.820 1.380 2.100 ;
        RECT  2.140 1.070 2.300 2.100 ;
        RECT  1.180 1.940 2.300 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.400 2.400 ;
        RECT  3.890 1.110 7.600 2.400 ;
        RECT  0.000 1.260 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.110 ;
        RECT  0.000 0.000 3.890 1.140 ;
        RECT  0.400 0.000 3.890 1.260 ;
    END
END BUFTM12HM

MACRO BUFM8HM
    CLASS CORE ;
    FOREIGN BUFM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.935  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.060 0.300 1.260 ;
        LAYER ME2 ;
        RECT  0.100 0.840 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.100 0.980 0.580 1.340 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 0.390 2.420 2.080 ;
        RECT  1.180 1.440 2.420 1.640 ;
        RECT  2.100 0.660 2.420 1.640 ;
        RECT  1.180 0.660 2.420 0.860 ;
        RECT  1.180 1.440 1.380 2.080 ;
        RECT  1.180 0.390 1.380 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.740 1.470 2.940 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.740 -0.140 2.940 0.660 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.310 0.340 0.820 ;
        RECT  0.140 0.660 0.960 0.820 ;
        RECT  0.760 1.040 1.760 1.240 ;
        RECT  0.760 0.660 0.960 1.720 ;
        RECT  0.140 1.520 0.960 1.720 ;
        RECT  0.140 1.520 0.340 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END BUFM8HM

MACRO BUFM6HM
    CLASS CORE ;
    FOREIGN BUFM6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.040  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.100 0.700 1.300 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.250 1.040 0.800 1.360 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.390 2.700 2.090 ;
        RECT  1.420 1.440 2.700 1.640 ;
        RECT  1.420 0.660 2.700 0.860 ;
        RECT  1.420 1.440 1.620 2.080 ;
        RECT  1.420 0.390 1.620 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.940 1.840 2.140 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        RECT  0.860 -0.140 1.140 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 0.380 0.580 0.860 ;
        RECT  0.380 0.680 1.200 0.860 ;
        RECT  1.000 1.040 2.300 1.240 ;
        RECT  1.000 0.680 1.200 1.740 ;
        RECT  0.340 1.540 1.200 1.740 ;
        RECT  0.340 1.540 0.630 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END BUFM6HM

MACRO BUFM5HM
    CLASS CORE ;
    FOREIGN BUFM5HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.125  LAYER ME1  ;
        ANTENNAGATEAREA 0.125  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.625  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.100 0.700 1.300 ;
        LAYER ME2 ;
        RECT  0.500 0.840 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.250 1.040 0.800 1.360 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.773  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.350 2.700 1.960 ;
        RECT  1.420 1.540 2.700 1.740 ;
        RECT  1.420 0.660 2.700 0.860 ;
        RECT  1.420 1.540 1.620 1.960 ;
        RECT  1.420 0.350 1.620 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.500 ;
        RECT  0.860 -0.140 1.140 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.400 0.350 0.610 0.860 ;
        RECT  0.400 0.660 1.200 0.860 ;
        RECT  1.000 1.040 2.300 1.240 ;
        RECT  1.000 0.660 1.200 1.740 ;
        RECT  0.380 1.540 1.200 1.740 ;
        RECT  0.380 1.540 0.580 2.000 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END BUFM5HM

MACRO BUFM4HM
    CLASS CORE ;
    FOREIGN BUFM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 0.920 1.180 ;
        RECT  0.100 0.840 0.340 1.180 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 1.450 2.300 1.650 ;
        RECT  2.100 0.660 2.300 1.650 ;
        RECT  1.540 0.660 2.300 0.840 ;
        RECT  1.540 1.450 1.740 2.090 ;
        RECT  1.540 0.390 1.740 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  2.060 1.840 2.260 2.540 ;
        RECT  0.980 1.900 1.260 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  2.020 -0.140 2.300 0.500 ;
        RECT  0.980 -0.140 1.260 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.500 0.360 0.700 0.820 ;
        RECT  0.500 0.660 1.350 0.820 ;
        RECT  1.170 1.010 1.900 1.290 ;
        RECT  1.170 0.660 1.350 1.740 ;
        RECT  0.500 1.580 1.350 1.740 ;
        RECT  0.500 1.580 0.700 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END BUFM4HM

MACRO BUFM48HM
    CLASS CORE ;
    FOREIGN BUFM48HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.893  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 3.150 1.220 ;
        RECT  0.100 0.760 0.410 1.220 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.878  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  15.160 1.500 15.460 2.080 ;
        RECT  3.780 0.660 15.420 0.860 ;
        RECT  15.220 0.330 15.420 0.860 ;
        RECT  3.740 1.500 15.460 1.740 ;
        RECT  14.180 1.500 14.380 2.080 ;
        RECT  14.180 0.320 14.380 0.860 ;
        RECT  13.140 1.500 13.340 2.080 ;
        RECT  13.140 0.390 13.340 0.860 ;
        RECT  12.100 1.500 12.300 2.080 ;
        RECT  12.100 0.390 12.300 0.860 ;
        RECT  11.060 1.500 11.260 2.080 ;
        RECT  11.060 0.390 11.260 0.860 ;
        RECT  10.020 1.500 10.220 2.080 ;
        RECT  10.020 0.390 10.220 0.860 ;
        RECT  9.650 0.660 9.950 1.740 ;
        RECT  8.980 1.500 9.180 2.080 ;
        RECT  8.980 0.390 9.180 0.860 ;
        RECT  7.940 1.500 8.140 2.080 ;
        RECT  7.940 0.390 8.140 0.860 ;
        RECT  6.900 1.500 7.100 2.080 ;
        RECT  6.900 0.390 7.100 0.860 ;
        RECT  5.860 1.500 6.060 2.080 ;
        RECT  5.860 0.390 6.060 0.860 ;
        RECT  4.820 1.500 5.020 2.080 ;
        RECT  4.820 0.390 5.020 0.860 ;
        RECT  3.740 1.500 3.980 2.080 ;
        RECT  3.780 0.390 3.980 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 15.600 2.540 ;
        RECT  14.660 1.900 14.940 2.540 ;
        RECT  13.620 1.900 13.900 2.540 ;
        RECT  12.580 1.900 12.860 2.540 ;
        RECT  11.540 1.900 11.820 2.540 ;
        RECT  10.500 1.900 10.780 2.540 ;
        RECT  9.460 1.900 9.740 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 15.600 0.140 ;
        RECT  14.660 -0.140 14.940 0.500 ;
        RECT  13.620 -0.140 13.900 0.500 ;
        RECT  12.580 -0.140 12.860 0.500 ;
        RECT  11.540 -0.140 11.820 0.500 ;
        RECT  10.500 -0.140 10.780 0.500 ;
        RECT  9.460 -0.140 9.740 0.500 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.100 -0.140 0.380 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.390 0.860 0.860 ;
        RECT  1.700 0.390 1.900 0.860 ;
        RECT  2.740 0.390 2.940 0.860 ;
        RECT  0.660 0.660 3.560 0.860 ;
        RECT  3.360 1.020 9.260 1.220 ;
        RECT  3.360 0.660 3.560 1.740 ;
        RECT  0.620 1.500 3.560 1.740 ;
        RECT  0.620 1.500 0.860 2.080 ;
        RECT  1.700 1.500 1.900 2.080 ;
        RECT  2.740 1.500 2.940 2.080 ;
        RECT  10.260 1.020 14.950 1.220 ;
        LAYER VTPH ;
        RECT  0.000 1.140 15.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 15.600 1.140 ;
    END
END BUFM48HM

MACRO BUFM40HM
    CLASS CORE ;
    FOREIGN BUFM40HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.744  LAYER ME2  ;
        ANTENNAGATEAREA 0.744  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.719  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.750 1.500 1.380 ;
        LAYER ME1 ;
        RECT  0.500 0.980 2.660 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.886  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  12.580 1.540 12.860 2.080 ;
        RECT  3.260 0.660 12.820 0.820 ;
        RECT  12.620 0.300 12.820 0.820 ;
        RECT  3.220 1.540 12.860 1.740 ;
        RECT  11.540 1.540 11.820 2.100 ;
        RECT  11.580 0.390 11.780 0.820 ;
        RECT  10.500 1.540 10.780 2.100 ;
        RECT  10.540 0.390 10.740 0.820 ;
        RECT  9.460 1.540 9.740 2.100 ;
        RECT  9.500 0.390 9.700 0.820 ;
        RECT  8.420 1.540 8.700 2.100 ;
        RECT  8.460 0.390 8.660 0.820 ;
        RECT  8.050 0.660 8.350 1.740 ;
        RECT  7.380 1.540 7.660 2.100 ;
        RECT  7.420 0.390 7.620 0.820 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  6.380 0.390 6.580 0.820 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.390 5.540 0.820 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.390 4.500 0.820 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  3.260 0.390 3.460 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  12.060 1.900 12.340 2.540 ;
        RECT  11.020 1.900 11.300 2.540 ;
        RECT  9.980 1.900 10.260 2.540 ;
        RECT  8.940 1.900 9.220 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.840 2.980 2.540 ;
        RECT  1.660 1.840 1.940 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  12.060 -0.140 12.340 0.500 ;
        RECT  11.020 -0.140 11.300 0.500 ;
        RECT  9.980 -0.140 10.260 0.500 ;
        RECT  8.940 -0.140 9.220 0.500 ;
        RECT  7.900 -0.140 8.180 0.500 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  2.220 0.380 2.420 0.820 ;
        RECT  0.140 0.660 3.040 0.820 ;
        RECT  2.840 0.980 7.660 1.180 ;
        RECT  2.840 0.660 3.040 1.680 ;
        RECT  0.100 1.480 3.040 1.680 ;
        RECT  0.100 1.480 0.380 2.100 ;
        RECT  1.140 1.480 1.420 2.100 ;
        RECT  2.180 1.480 2.460 2.100 ;
        RECT  8.660 0.980 12.180 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.140 ;
    END
END BUFM40HM

MACRO BUFM3HM
    CLASS CORE ;
    FOREIGN BUFM3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.271  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.380 1.020 0.580 1.220 ;
        LAYER ME2 ;
        RECT  0.380 0.750 0.700 1.380 ;
        LAYER ME1 ;
        RECT  0.300 0.980 0.660 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.377  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 1.540 2.300 1.740 ;
        RECT  2.100 0.660 2.300 1.740 ;
        RECT  1.280 0.660 2.300 0.820 ;
        RECT  1.280 1.540 1.480 2.020 ;
        RECT  1.280 0.390 1.480 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.760 1.900 2.040 2.540 ;
        RECT  0.760 1.840 0.960 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.760 -0.140 2.040 0.500 ;
        RECT  0.720 -0.140 1.000 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.240 0.300 0.440 0.820 ;
        RECT  0.240 0.660 1.060 0.820 ;
        RECT  0.860 1.060 1.700 1.260 ;
        RECT  0.860 0.660 1.060 1.680 ;
        RECT  0.240 1.480 1.060 1.680 ;
        RECT  0.240 1.480 0.440 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END BUFM3HM

MACRO BUFM36HM
    CLASS CORE ;
    FOREIGN BUFM36HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.744  LAYER ME2  ;
        ANTENNAGATEAREA 0.744  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.950  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.750 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.150 0.980 2.640 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.464  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.540 1.540 11.820 2.100 ;
        RECT  3.260 0.660 11.780 0.820 ;
        RECT  11.580 0.390 11.780 0.820 ;
        RECT  3.220 1.540 11.820 1.740 ;
        RECT  10.500 1.540 10.780 2.100 ;
        RECT  10.540 0.390 10.740 0.820 ;
        RECT  9.460 1.540 9.740 2.100 ;
        RECT  9.500 0.390 9.700 0.820 ;
        RECT  8.420 1.540 8.700 2.100 ;
        RECT  8.460 0.390 8.660 0.820 ;
        RECT  8.050 0.660 8.350 1.740 ;
        RECT  7.380 1.540 7.660 2.100 ;
        RECT  7.420 0.390 7.620 0.820 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  6.380 0.390 6.580 0.820 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.390 5.540 0.820 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.390 4.500 0.820 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  3.260 0.390 3.460 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 12.800 2.540 ;
        RECT  12.100 1.480 12.300 2.540 ;
        RECT  11.020 1.900 11.300 2.540 ;
        RECT  9.980 1.900 10.260 2.540 ;
        RECT  8.940 1.900 9.220 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.840 2.980 2.540 ;
        RECT  1.660 1.840 1.940 2.540 ;
        RECT  0.620 1.840 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 12.800 0.140 ;
        RECT  12.060 -0.140 12.340 0.580 ;
        RECT  11.020 -0.140 11.300 0.500 ;
        RECT  9.980 -0.140 10.260 0.500 ;
        RECT  8.940 -0.140 9.220 0.500 ;
        RECT  7.900 -0.140 8.180 0.500 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  2.220 0.380 2.420 0.820 ;
        RECT  0.140 0.660 3.040 0.820 ;
        RECT  2.840 0.980 7.660 1.180 ;
        RECT  2.840 0.660 3.040 1.680 ;
        RECT  0.100 1.480 3.040 1.680 ;
        RECT  0.100 1.480 0.380 2.100 ;
        RECT  1.140 1.480 1.420 2.100 ;
        RECT  2.180 1.480 2.460 2.100 ;
        RECT  8.660 0.980 11.950 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 12.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 12.800 1.140 ;
    END
END BUFM36HM

MACRO BUFM32HM
    CLASS CORE ;
    FOREIGN BUFM32HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.394  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.750 1.500 1.380 ;
        LAYER ME1 ;
        RECT  0.200 0.980 2.640 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.968  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.500 1.540 10.780 2.100 ;
        RECT  3.260 0.660 10.740 0.820 ;
        RECT  10.540 0.390 10.740 0.820 ;
        RECT  3.220 1.540 10.780 1.740 ;
        RECT  9.460 1.540 9.740 2.100 ;
        RECT  9.500 0.390 9.700 0.820 ;
        RECT  8.420 1.540 8.700 2.100 ;
        RECT  8.460 0.390 8.660 0.820 ;
        RECT  8.050 0.660 8.350 1.740 ;
        RECT  7.380 1.540 7.660 2.100 ;
        RECT  7.420 0.390 7.620 0.820 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  6.380 0.390 6.580 0.820 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.390 5.540 0.820 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.390 4.500 0.820 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  3.260 0.390 3.460 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  11.060 1.480 11.260 2.540 ;
        RECT  9.980 1.900 10.260 2.540 ;
        RECT  8.940 1.900 9.220 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.740 1.840 2.940 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.060 -0.140 11.260 0.670 ;
        RECT  9.980 -0.140 10.260 0.500 ;
        RECT  8.940 -0.140 9.220 0.500 ;
        RECT  7.900 -0.140 8.180 0.500 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  2.220 0.380 2.420 0.820 ;
        RECT  0.140 0.660 3.040 0.820 ;
        RECT  2.840 0.980 7.660 1.180 ;
        RECT  2.840 0.660 3.040 1.680 ;
        RECT  0.140 1.480 3.040 1.680 ;
        RECT  0.140 1.480 0.340 2.000 ;
        RECT  1.180 1.480 1.380 2.000 ;
        RECT  2.220 1.480 2.420 2.000 ;
        RECT  8.660 0.980 10.890 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.140 ;
    END
END BUFM32HM

MACRO BUFM2HM
    CLASS CORE ;
    FOREIGN BUFM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.899  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.040 0.300 1.240 ;
        LAYER ME2 ;
        RECT  0.100 0.750 0.300 1.380 ;
        LAYER ME1 ;
        RECT  0.100 0.980 0.560 1.300 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.140 1.800 1.500 2.000 ;
        RECT  1.300 0.350 1.500 2.000 ;
        RECT  1.140 0.350 1.500 0.550 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 1.600 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 1.600 0.140 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.300 0.340 0.820 ;
        RECT  0.140 0.660 1.020 0.820 ;
        RECT  0.860 0.660 1.020 1.680 ;
        RECT  0.140 1.480 1.020 1.680 ;
        RECT  0.140 1.480 0.340 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 1.600 1.140 ;
    END
END BUFM2HM

MACRO BUFM28HM
    CLASS CORE ;
    FOREIGN BUFM28HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.782  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.750 1.500 1.380 ;
        LAYER ME1 ;
        RECT  0.380 0.980 2.120 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.472  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.940 1.540 9.220 2.100 ;
        RECT  2.740 0.660 9.180 0.820 ;
        RECT  8.980 0.390 9.180 0.820 ;
        RECT  2.700 1.540 9.220 1.740 ;
        RECT  7.900 1.540 8.180 2.100 ;
        RECT  7.940 0.390 8.140 0.820 ;
        RECT  7.600 0.660 7.920 1.740 ;
        RECT  6.860 1.540 7.140 2.100 ;
        RECT  6.900 0.390 7.100 0.820 ;
        RECT  5.820 1.540 6.100 2.100 ;
        RECT  5.860 0.390 6.060 0.820 ;
        RECT  4.780 1.540 5.060 2.100 ;
        RECT  4.820 0.390 5.020 0.820 ;
        RECT  3.740 1.540 4.020 2.100 ;
        RECT  3.780 0.390 3.980 0.820 ;
        RECT  2.700 1.540 2.980 2.100 ;
        RECT  2.740 0.390 2.940 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.500 1.480 9.700 2.540 ;
        RECT  8.420 1.900 8.700 2.540 ;
        RECT  7.380 1.900 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.220 1.840 2.420 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.500 -0.140 9.700 0.660 ;
        RECT  8.420 -0.140 8.700 0.500 ;
        RECT  7.380 -0.140 7.660 0.500 ;
        RECT  6.340 -0.140 6.620 0.500 ;
        RECT  5.300 -0.140 5.580 0.500 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.380 0.860 0.820 ;
        RECT  1.700 0.380 1.900 0.820 ;
        RECT  0.660 0.660 2.520 0.820 ;
        RECT  2.320 0.980 7.140 1.180 ;
        RECT  2.320 0.660 2.520 1.660 ;
        RECT  0.660 1.460 2.520 1.660 ;
        RECT  0.660 1.460 0.860 2.100 ;
        RECT  1.700 1.460 1.900 2.100 ;
        RECT  8.140 0.980 9.280 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
    END
END BUFM28HM

MACRO BUFM24HM
    CLASS CORE ;
    FOREIGN BUFM24HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.957  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.750 1.100 1.380 ;
        LAYER ME1 ;
        RECT  0.220 0.980 1.600 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.976  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.380 0.390 7.660 2.100 ;
        RECT  2.180 1.540 7.660 1.740 ;
        RECT  7.130 0.660 7.660 1.740 ;
        RECT  2.220 0.660 7.660 0.820 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  6.380 0.390 6.580 0.820 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.390 5.540 0.820 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.390 4.500 0.820 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  3.260 0.390 3.460 0.820 ;
        RECT  2.180 1.540 2.460 2.100 ;
        RECT  2.220 0.390 2.420 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.940 1.480 8.140 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.940 -0.140 8.140 0.660 ;
        RECT  6.860 -0.140 7.140 0.500 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  0.140 0.660 2.000 0.820 ;
        RECT  1.800 0.980 6.620 1.180 ;
        RECT  0.140 1.460 2.000 1.660 ;
        RECT  1.800 0.660 2.000 1.680 ;
        RECT  1.180 1.460 2.000 1.680 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.180 1.460 1.380 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END BUFM24HM

MACRO BUFM20HM
    CLASS CORE ;
    FOREIGN BUFM20HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.934  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.750 1.100 1.380 ;
        LAYER ME1 ;
        RECT  0.240 0.980 1.600 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.480  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  2.220 0.660 6.580 0.820 ;
        RECT  6.380 0.390 6.580 0.820 ;
        RECT  2.180 1.540 6.620 1.740 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.390 5.540 0.820 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.390 4.500 0.820 ;
        RECT  4.050 0.660 4.350 1.740 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  3.260 0.390 3.460 0.820 ;
        RECT  2.180 1.540 2.460 2.100 ;
        RECT  2.220 0.390 2.420 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  6.900 1.480 7.100 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.900 -0.140 7.100 0.660 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  0.140 0.660 2.000 0.820 ;
        RECT  1.800 0.980 3.830 1.180 ;
        RECT  1.800 0.660 2.000 1.660 ;
        RECT  0.140 1.460 2.000 1.660 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  1.180 1.460 1.380 2.100 ;
        RECT  4.960 0.980 6.700 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END BUFM20HM

MACRO BUFM18HM
    CLASS CORE ;
    FOREIGN BUFM18HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.446  LAYER ME2  ;
        ANTENNAGATEAREA 0.446  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.689  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.750 1.100 1.380 ;
        LAYER ME1 ;
        RECT  0.450 0.980 1.600 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.406  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 1.540 6.620 2.100 ;
        RECT  2.220 0.660 6.620 0.820 ;
        RECT  6.340 0.390 6.620 0.820 ;
        RECT  2.180 1.540 6.620 1.740 ;
        RECT  5.300 1.540 5.580 2.100 ;
        RECT  5.340 0.390 5.540 0.820 ;
        RECT  4.260 1.540 4.540 2.100 ;
        RECT  4.300 0.390 4.500 0.820 ;
        RECT  4.050 0.660 4.350 1.740 ;
        RECT  3.220 1.540 3.500 2.100 ;
        RECT  3.260 0.390 3.460 0.820 ;
        RECT  2.180 1.540 2.460 2.100 ;
        RECT  2.220 0.390 2.420 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.700 1.840 1.900 2.540 ;
        RECT  0.660 1.840 0.860 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.820 -0.140 6.100 0.500 ;
        RECT  4.780 -0.140 5.060 0.500 ;
        RECT  3.740 -0.140 4.020 0.500 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.660 -0.140 1.940 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 0.340 0.820 ;
        RECT  1.180 0.380 1.380 0.820 ;
        RECT  0.140 0.660 2.000 0.820 ;
        RECT  1.800 0.980 3.780 1.180 ;
        RECT  0.140 1.460 2.000 1.660 ;
        RECT  1.800 0.660 2.000 1.680 ;
        RECT  1.180 1.460 2.000 1.680 ;
        RECT  1.180 1.460 1.380 2.080 ;
        RECT  0.140 1.460 0.340 2.100 ;
        RECT  4.610 0.980 6.250 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END BUFM18HM

MACRO BUFM16HM
    CLASS CORE ;
    FOREIGN BUFM16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.642  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.020 0.700 1.220 ;
        LAYER ME2 ;
        RECT  0.500 0.750 0.700 1.380 ;
        LAYER ME1 ;
        RECT  0.440 0.980 1.080 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.780 1.540 5.060 2.100 ;
        RECT  1.700 0.660 5.060 0.820 ;
        RECT  4.780 0.390 5.060 0.820 ;
        RECT  1.660 1.540 5.060 1.740 ;
        RECT  3.740 1.540 4.020 2.100 ;
        RECT  3.780 0.390 3.980 0.820 ;
        RECT  3.650 0.660 3.900 1.740 ;
        RECT  2.700 1.540 2.980 2.100 ;
        RECT  2.740 0.390 2.940 0.820 ;
        RECT  1.660 1.540 1.940 2.100 ;
        RECT  1.700 0.390 1.900 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.340 1.480 5.540 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.340 -0.140 5.540 0.670 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.380 0.860 0.820 ;
        RECT  0.660 0.660 1.480 0.820 ;
        RECT  1.280 0.980 3.260 1.180 ;
        RECT  1.280 0.660 1.480 1.660 ;
        RECT  0.660 1.460 1.480 1.660 ;
        RECT  0.660 1.460 0.860 2.100 ;
        RECT  4.120 0.980 5.240 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END BUFM16HM

MACRO BUFM14HM
    CLASS CORE ;
    FOREIGN BUFM14HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 1.080 1.180 ;
        RECT  0.100 0.790 0.390 1.180 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.910  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.780 1.540 5.060 2.100 ;
        RECT  1.700 0.660 5.060 0.820 ;
        RECT  4.780 0.390 5.060 0.820 ;
        RECT  1.660 1.540 5.060 1.740 ;
        RECT  3.740 1.540 4.020 2.100 ;
        RECT  3.780 0.390 3.980 0.820 ;
        RECT  3.250 0.660 3.550 1.740 ;
        RECT  2.700 1.540 2.980 2.100 ;
        RECT  2.740 0.390 2.940 0.820 ;
        RECT  1.660 1.540 1.940 2.100 ;
        RECT  1.700 0.390 1.900 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.180 1.840 1.380 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.260 -0.140 4.540 0.500 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.380 0.860 0.820 ;
        RECT  0.660 0.660 1.480 0.820 ;
        RECT  1.280 0.980 2.860 1.180 ;
        RECT  1.280 0.660 1.480 1.680 ;
        RECT  0.660 1.460 1.480 1.680 ;
        RECT  0.660 1.460 0.860 2.100 ;
        RECT  4.000 0.980 4.720 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END BUFM14HM

MACRO BUFM12HM
    CLASS CORE ;
    FOREIGN BUFM12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.747  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.750 1.100 1.380 ;
        LAYER ME1 ;
        RECT  0.480 0.980 1.180 1.280 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.840 1.540 4.120 2.100 ;
        RECT  1.800 0.660 4.080 0.820 ;
        RECT  3.880 0.390 4.080 0.820 ;
        RECT  1.760 1.540 4.120 1.740 ;
        RECT  2.800 1.540 3.080 2.100 ;
        RECT  2.840 0.390 3.040 0.820 ;
        RECT  2.430 0.660 2.790 1.740 ;
        RECT  1.760 1.540 2.040 2.100 ;
        RECT  1.800 0.390 2.000 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.400 1.480 4.600 2.540 ;
        RECT  3.320 1.900 3.600 2.540 ;
        RECT  2.280 1.900 2.560 2.540 ;
        RECT  1.280 1.840 1.480 2.540 ;
        RECT  0.240 1.480 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.400 -0.140 4.600 0.670 ;
        RECT  3.320 -0.140 3.600 0.500 ;
        RECT  2.280 -0.140 2.560 0.500 ;
        RECT  1.240 -0.140 1.520 0.500 ;
        RECT  0.240 -0.140 0.440 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.760 0.380 0.960 0.820 ;
        RECT  0.760 0.660 1.580 0.820 ;
        RECT  1.380 0.980 2.270 1.180 ;
        RECT  1.380 0.660 1.580 1.660 ;
        RECT  0.760 1.460 1.580 1.660 ;
        RECT  0.760 1.460 0.960 2.100 ;
        RECT  3.220 0.980 4.300 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END BUFM12HM

MACRO BUFM10HM
    CLASS CORE ;
    FOREIGN BUFM10HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.414  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.840 1.540 4.120 2.100 ;
        RECT  1.800 0.660 4.080 0.820 ;
        RECT  3.880 0.390 4.080 0.820 ;
        RECT  1.760 1.540 4.120 1.740 ;
        RECT  2.800 1.540 3.080 2.100 ;
        RECT  2.840 0.390 3.040 0.820 ;
        RECT  2.500 0.660 2.700 1.740 ;
        RECT  1.760 1.540 2.040 2.100 ;
        RECT  1.800 0.390 2.000 0.820 ;
        END
    END Z
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.251  LAYER ME1  ;
        ANTENNAGATEAREA 0.251  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.073  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.750 1.100 1.380 ;
        LAYER ME1 ;
        RECT  0.480 0.980 1.180 1.280 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.320 1.900 3.600 2.540 ;
        RECT  2.280 1.900 2.560 2.540 ;
        RECT  1.280 1.840 1.480 2.540 ;
        RECT  0.240 1.680 0.440 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.320 -0.140 3.600 0.500 ;
        RECT  2.280 -0.140 2.560 0.500 ;
        RECT  1.240 -0.140 1.520 0.500 ;
        RECT  0.200 -0.140 0.480 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.720 0.380 1.000 0.820 ;
        RECT  0.720 0.660 1.580 0.820 ;
        RECT  1.380 0.980 2.270 1.180 ;
        RECT  1.380 0.660 1.580 1.680 ;
        RECT  0.760 1.480 1.580 1.680 ;
        RECT  0.760 1.480 0.960 1.960 ;
        RECT  3.010 0.980 3.750 1.180 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END BUFM10HM

MACRO BHDM1HM
    CLASS CORE ;
    FOREIGN BHDM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.189  LAYER ME1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.053  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.520 1.680 1.900 1.840 ;
        RECT  1.680 0.560 1.900 1.840 ;
        RECT  0.520 1.080 0.720 1.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  0.740 2.020 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  0.740 -0.140 0.940 0.460 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.620 1.400 0.820 ;
        RECT  1.200 0.620 1.400 1.360 ;
        RECT  0.100 0.620 0.340 1.900 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END BHDM1HM

MACRO AOI33M8HM
    CLASS CORE ;
    FOREIGN AOI33M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.223  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  8.100 1.020 8.300 1.220 ;
        LAYER ME2 ;
        RECT  8.100 0.770 8.300 1.470 ;
        LAYER ME1 ;
        RECT  7.500 0.980 8.580 1.300 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.020 5.900 1.220 ;
        LAYER ME2 ;
        RECT  5.700 0.770 5.900 1.470 ;
        LAYER ME1 ;
        RECT  4.760 0.980 6.240 1.300 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.080 1.260 12.740 1.420 ;
        RECT  12.460 0.840 12.740 1.420 ;
        RECT  10.760 1.120 11.040 1.420 ;
        RECT  9.080 1.020 9.240 1.420 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.581  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.520 0.800 11.800 1.100 ;
        RECT  9.600 0.800 11.800 0.960 ;
        RECT  9.600 0.800 9.960 1.100 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.600 1.260 4.320 1.420 ;
        RECT  4.060 0.840 4.320 1.420 ;
        RECT  2.360 1.120 2.640 1.420 ;
        RECT  0.600 1.000 0.910 1.420 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.581  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.120 0.800 3.400 1.100 ;
        RECT  1.200 0.800 3.400 0.960 ;
        RECT  1.200 0.800 1.560 1.100 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.528  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.990 1.580 12.620 1.740 ;
        RECT  4.740 0.660 8.620 0.820 ;
        RECT  8.340 0.620 8.620 0.820 ;
        RECT  7.300 0.620 7.580 0.820 ;
        RECT  6.990 0.660 7.160 1.740 ;
        RECT  6.840 0.660 7.160 1.100 ;
        RECT  5.780 0.620 6.060 0.820 ;
        RECT  4.740 0.620 5.020 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.200 2.540 ;
        RECT  5.980 1.900 6.260 2.540 ;
        RECT  4.940 1.900 5.220 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        RECT  1.820 1.900 2.100 2.540 ;
        RECT  0.780 1.900 1.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.200 0.140 ;
        RECT  11.740 -0.140 12.020 0.320 ;
        RECT  9.860 -0.140 10.140 0.320 ;
        RECT  3.340 -0.140 3.620 0.320 ;
        RECT  1.460 -0.140 1.740 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.260 0.300 6.580 0.460 ;
        RECT  5.260 0.300 5.540 0.500 ;
        RECT  6.300 0.300 6.580 0.500 ;
        RECT  4.260 0.300 4.460 0.640 ;
        RECT  0.420 0.480 4.460 0.640 ;
        RECT  6.780 0.300 9.160 0.460 ;
        RECT  8.860 0.300 9.160 0.640 ;
        RECT  6.780 0.300 7.060 0.500 ;
        RECT  7.820 0.300 8.100 0.500 ;
        RECT  8.860 0.480 12.940 0.640 ;
        RECT  0.220 1.580 6.800 1.740 ;
        RECT  6.560 1.580 6.800 2.060 ;
        RECT  12.860 1.730 13.060 2.060 ;
        RECT  6.560 1.900 13.060 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 13.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.200 1.140 ;
    END
END AOI33M8HM

MACRO AOI33M4HM
    CLASS CORE ;
    FOREIGN AOI33M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.642  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.130 5.500 1.330 ;
        LAYER ME2 ;
        RECT  5.300 0.820 5.500 1.500 ;
        LAYER ME1 ;
        RECT  5.160 1.120 5.880 1.340 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.817  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.060 2.700 1.260 ;
        LAYER ME2 ;
        RECT  2.500 0.820 2.700 1.440 ;
        LAYER ME1 ;
        RECT  2.390 1.000 3.100 1.330 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.136  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.060 3.900 1.260 ;
        LAYER ME2 ;
        RECT  3.700 0.820 3.900 1.440 ;
        LAYER ME1 ;
        RECT  3.620 1.000 3.940 1.330 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.100 0.800 6.360 1.280 ;
        RECT  4.740 0.800 6.360 0.960 ;
        RECT  4.740 0.800 4.940 1.280 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.800 0.800 2.050 1.260 ;
        RECT  0.400 0.800 2.050 0.960 ;
        RECT  0.400 0.800 0.700 1.360 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.264  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.780 1.580 6.220 1.740 ;
        RECT  4.100 0.620 4.300 1.740 ;
        RECT  2.490 0.660 4.300 0.820 ;
        RECT  4.020 0.620 4.300 0.820 ;
        RECT  2.490 0.620 2.780 0.820 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.642  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 0.820 1.500 1.440 ;
        LAYER ME1 ;
        RECT  0.880 1.120 1.600 1.340 ;
        END
    END B3
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  5.420 -0.140 5.700 0.320 ;
        RECT  1.100 -0.140 1.380 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.020 0.300 3.300 0.460 ;
        RECT  3.020 0.300 3.300 0.500 ;
        RECT  2.020 0.300 2.220 0.640 ;
        RECT  0.180 0.480 2.220 0.640 ;
        RECT  3.500 0.300 4.780 0.460 ;
        RECT  4.570 0.300 4.780 0.640 ;
        RECT  3.500 0.300 3.800 0.500 ;
        RECT  4.570 0.480 6.620 0.640 ;
        RECT  0.140 1.580 3.500 1.740 ;
        RECT  3.300 1.580 3.500 2.060 ;
        RECT  0.140 1.580 0.340 1.910 ;
        RECT  6.460 1.690 6.660 2.060 ;
        RECT  3.300 1.900 6.660 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END AOI33M4HM

MACRO AOI33M2HM
    CLASS CORE ;
    FOREIGN AOI33M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.810 1.600 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.820 1.120 1.260 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.820 0.700 1.260 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.000 0.840 2.300 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.800 2.700 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.810 3.140 1.300 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.862  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 1.500 3.500 2.100 ;
        RECT  3.300 0.480 3.500 2.100 ;
        RECT  1.660 0.480 3.500 0.640 ;
        RECT  2.140 1.500 3.500 1.660 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.180 -0.140 3.460 0.320 ;
        RECT  0.260 -0.140 0.460 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 1.520 1.940 1.740 ;
        RECT  1.650 1.520 1.940 2.100 ;
        RECT  0.620 1.520 0.900 2.100 ;
        RECT  2.700 1.820 2.980 2.100 ;
        RECT  1.650 1.940 2.980 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI33M2HM

MACRO AOI33M1HM
    CLASS CORE ;
    FOREIGN AOI33M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.810 1.640 1.290 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.820 1.120 1.340 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.370 0.820 0.700 1.340 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.880 0.840 2.300 1.300 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.800 2.700 1.300 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.810 3.140 1.300 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.611  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 1.470 3.500 1.960 ;
        RECT  3.300 0.480 3.500 1.960 ;
        RECT  2.860 0.480 3.500 0.640 ;
        RECT  2.180 1.470 3.500 1.660 ;
        RECT  1.660 0.340 3.020 0.500 ;
        RECT  2.180 1.470 2.460 1.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.740 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.180 -0.140 3.460 0.320 ;
        RECT  0.260 -0.140 0.460 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.520 1.900 1.740 ;
        RECT  1.700 1.520 1.900 2.100 ;
        RECT  0.660 1.520 0.860 2.020 ;
        RECT  2.700 1.820 2.980 2.100 ;
        RECT  1.700 1.940 2.980 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI33M1HM

MACRO AOI33M0HM
    CLASS CORE ;
    FOREIGN AOI33M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.810 1.640 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.880 0.820 1.120 1.260 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.370 0.820 0.700 1.260 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.880 0.840 2.300 1.240 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.800 2.700 1.240 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.810 3.140 1.240 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.486  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.400 3.500 1.940 ;
        RECT  3.300 0.480 3.500 1.940 ;
        RECT  2.860 0.480 3.500 0.640 ;
        RECT  2.180 1.400 3.500 1.560 ;
        RECT  1.660 0.340 3.020 0.500 ;
        RECT  2.180 1.400 2.460 1.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  1.140 1.820 1.420 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.180 -0.140 3.460 0.320 ;
        RECT  0.260 -0.140 0.460 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.490 1.900 1.660 ;
        RECT  1.700 1.490 1.900 2.100 ;
        RECT  0.660 1.490 0.860 2.010 ;
        RECT  2.700 1.720 2.980 2.100 ;
        RECT  1.700 1.940 2.980 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI33M0HM

MACRO AOI32M8HM
    CLASS CORE ;
    FOREIGN AOI32M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.020 5.900 1.220 ;
        LAYER ME2 ;
        RECT  5.700 0.780 5.900 1.500 ;
        LAYER ME1 ;
        RECT  4.840 0.980 6.320 1.300 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.080 1.260 10.740 1.420 ;
        RECT  10.460 0.840 10.740 1.420 ;
        RECT  8.760 1.120 9.040 1.420 ;
        RECT  7.080 1.020 7.240 1.420 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.581  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.520 0.800 9.860 1.100 ;
        RECT  7.600 0.800 9.860 0.960 ;
        RECT  7.600 0.800 7.960 1.100 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.260 4.320 1.420 ;
        RECT  4.060 0.840 4.320 1.420 ;
        RECT  2.360 1.120 2.640 1.420 ;
        RECT  0.660 1.060 0.860 1.420 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.120 0.800 3.400 1.100 ;
        RECT  1.200 0.800 3.400 0.960 ;
        RECT  1.200 0.800 1.560 1.100 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.698  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.980 1.580 10.620 1.740 ;
        RECT  6.500 0.620 6.700 1.740 ;
        RECT  4.500 0.660 6.700 0.820 ;
        RECT  6.380 0.620 6.700 0.820 ;
        RECT  5.340 0.620 5.620 0.820 ;
        RECT  4.500 0.480 4.660 0.820 ;
        RECT  0.420 0.480 4.660 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        RECT  1.820 1.900 2.100 2.540 ;
        RECT  0.780 1.900 1.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  9.740 -0.140 10.020 0.320 ;
        RECT  7.860 -0.140 8.140 0.320 ;
        RECT  3.340 -0.140 3.620 0.320 ;
        RECT  1.460 -0.140 1.740 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  4.820 0.300 7.160 0.460 ;
        RECT  6.860 0.300 7.160 0.640 ;
        RECT  4.820 0.300 5.100 0.500 ;
        RECT  5.860 0.300 6.140 0.500 ;
        RECT  6.860 0.480 10.940 0.640 ;
        RECT  0.220 1.580 4.780 1.740 ;
        RECT  4.500 1.580 4.780 2.060 ;
        RECT  10.860 1.730 11.060 2.060 ;
        RECT  4.500 1.900 11.060 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
    END
END AOI32M8HM

MACRO AOI32M4HM
    CLASS CORE ;
    FOREIGN AOI32M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.690  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 0.820 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.880 1.120 1.600 1.340 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.468  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.060 2.700 1.260 ;
        LAYER ME2 ;
        RECT  2.500 0.820 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.300 1.000 2.810 1.330 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.760 1.260 5.540 1.420 ;
        RECT  5.240 0.840 5.540 1.420 ;
        RECT  3.760 1.020 3.920 1.420 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.290  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.280 0.800 4.810 1.100 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.840 0.800 2.040 1.220 ;
        RECT  0.400 0.800 2.040 0.960 ;
        RECT  0.400 0.800 0.700 1.340 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.555  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.580 5.420 1.740 ;
        RECT  3.030 1.240 3.560 1.740 ;
        RECT  3.030 0.680 3.380 1.740 ;
        RECT  3.060 0.620 3.380 1.740 ;
        RECT  2.210 0.680 3.380 0.840 ;
        RECT  2.210 0.480 2.370 0.840 ;
        RECT  0.180 0.480 2.370 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  4.540 -0.140 4.820 0.320 ;
        RECT  1.100 -0.140 1.380 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.530 0.300 3.780 0.460 ;
        RECT  3.580 0.300 3.780 0.640 ;
        RECT  2.530 0.300 2.820 0.500 ;
        RECT  3.580 0.480 5.740 0.640 ;
        RECT  0.140 1.580 2.460 1.740 ;
        RECT  2.180 1.580 2.460 2.060 ;
        RECT  0.140 1.580 0.340 1.960 ;
        RECT  5.660 1.640 5.860 2.060 ;
        RECT  2.180 1.900 5.860 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END AOI32M4HM

MACRO AOI32M2HM
    CLASS CORE ;
    FOREIGN AOI32M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.600 0.840 1.900 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.800 2.300 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.810 2.740 1.340 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.810 1.160 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.260 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.898  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 1.500 3.100 2.100 ;
        RECT  2.900 0.480 3.100 2.100 ;
        RECT  1.260 0.480 3.100 0.640 ;
        RECT  1.740 1.500 3.100 1.660 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  0.740 1.900 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.780 -0.140 3.060 0.320 ;
        RECT  0.260 -0.140 0.460 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 1.520 1.540 1.740 ;
        RECT  1.250 1.520 1.540 2.100 ;
        RECT  0.220 1.520 0.500 2.100 ;
        RECT  2.300 1.820 2.580 2.100 ;
        RECT  1.250 1.940 2.580 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AOI32M2HM

MACRO AOI32M1HM
    CLASS CORE ;
    FOREIGN AOI32M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.520 0.810 1.900 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.800 2.300 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.810 2.740 1.340 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.810 1.160 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.840 0.700 1.260 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.707  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.520 3.100 2.000 ;
        RECT  2.900 0.480 3.100 2.000 ;
        RECT  2.460 0.480 3.100 0.640 ;
        RECT  1.740 1.520 3.100 1.740 ;
        RECT  1.180 0.340 2.620 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.780 -0.140 3.060 0.320 ;
        RECT  0.180 -0.140 0.380 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 1.560 1.420 1.740 ;
        RECT  1.220 1.560 1.420 2.100 ;
        RECT  0.180 1.560 0.380 2.060 ;
        RECT  2.300 1.900 2.580 2.100 ;
        RECT  1.220 1.940 2.580 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AOI32M1HM

MACRO AOI32M0HM
    CLASS CORE ;
    FOREIGN AOI32M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.520 0.810 1.900 1.200 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.800 2.300 1.300 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.810 2.740 1.340 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.810 1.160 1.290 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 0.840 0.700 1.340 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 1.580 3.100 2.050 ;
        RECT  2.900 0.480 3.100 2.050 ;
        RECT  2.460 0.480 3.100 0.640 ;
        RECT  1.700 1.580 3.100 1.740 ;
        RECT  1.180 0.340 2.620 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  0.660 1.900 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.780 -0.140 3.060 0.320 ;
        RECT  0.180 -0.140 0.380 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 1.560 1.420 1.740 ;
        RECT  1.220 1.560 1.420 2.060 ;
        RECT  0.180 1.560 0.380 2.060 ;
        RECT  1.220 1.900 2.620 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AOI32M0HM

MACRO AOI31M8HM
    CLASS CORE ;
    FOREIGN AOI31M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        ANTENNAGATEAREA 0.595  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.573  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.700 1.020 3.900 1.220 ;
        LAYER ME2 ;
        RECT  3.700 0.780 3.900 1.500 ;
        LAYER ME1 ;
        RECT  2.840 0.980 4.320 1.300 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        ANTENNAGATEAREA 0.504  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.816  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.020 1.500 1.220 ;
        LAYER ME2 ;
        RECT  1.300 0.780 1.500 1.500 ;
        LAYER ME1 ;
        RECT  0.860 1.020 2.340 1.300 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.595  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.080 1.260 8.740 1.420 ;
        RECT  8.460 0.840 8.740 1.420 ;
        RECT  6.760 1.120 7.040 1.420 ;
        RECT  5.080 1.020 5.240 1.420 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.581  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.520 0.800 7.800 1.100 ;
        RECT  5.600 0.800 7.800 0.960 ;
        RECT  5.600 0.800 5.960 1.100 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.457  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.980 1.580 8.620 1.740 ;
        RECT  4.500 0.620 4.700 1.740 ;
        RECT  1.300 0.660 4.700 0.820 ;
        RECT  4.380 0.620 4.700 0.820 ;
        RECT  3.340 0.620 3.620 0.820 ;
        RECT  2.340 0.400 2.540 0.820 ;
        RECT  1.300 0.360 1.500 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.200 2.540 ;
        RECT  1.980 1.840 2.260 2.540 ;
        RECT  0.940 1.840 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.200 0.140 ;
        RECT  7.740 -0.140 8.020 0.320 ;
        RECT  5.860 -0.140 6.140 0.320 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        RECT  0.780 -0.140 0.980 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.820 0.300 5.160 0.460 ;
        RECT  4.860 0.300 5.160 0.640 ;
        RECT  2.820 0.300 3.100 0.500 ;
        RECT  3.860 0.300 4.140 0.500 ;
        RECT  4.860 0.480 8.940 0.640 ;
        RECT  0.420 1.470 2.780 1.660 ;
        RECT  2.500 1.470 2.780 2.060 ;
        RECT  8.860 1.800 9.100 2.060 ;
        RECT  2.500 1.900 9.100 2.060 ;
        RECT  0.420 1.470 0.700 2.100 ;
        RECT  1.460 1.470 1.740 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.200 1.140 ;
    END
END AOI31M8HM

MACRO AOI31M4HM
    CLASS CORE ;
    FOREIGN AOI31M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.625  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.020 1.900 1.220 ;
        LAYER ME2 ;
        RECT  1.700 0.810 1.900 1.400 ;
        LAYER ME1 ;
        RECT  1.560 1.020 2.200 1.310 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.747  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.020 3.500 1.220 ;
        LAYER ME2 ;
        RECT  3.300 0.810 3.500 1.400 ;
        LAYER ME1 ;
        RECT  3.080 0.980 3.720 1.340 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.850 1.020 5.100 1.560 ;
        RECT  4.120 1.020 5.100 1.220 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.740 1.540 4.580 1.740 ;
        RECT  2.360 1.200 2.700 1.740 ;
        RECT  2.360 0.620 2.580 1.740 ;
        RECT  0.220 0.660 2.580 0.820 ;
        RECT  2.260 0.620 2.580 0.820 ;
        RECT  1.260 0.310 1.460 0.820 ;
        RECT  0.220 0.310 0.420 0.820 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        ANTENNAGATEAREA 0.252  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.981  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.020 1.100 1.220 ;
        LAYER ME2 ;
        RECT  0.900 0.810 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.520 0.980 1.160 1.300 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.300 -0.140 4.580 0.500 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.740 0.300 3.540 0.460 ;
        RECT  1.740 0.300 2.020 0.500 ;
        RECT  3.260 0.300 3.540 0.500 ;
        RECT  2.740 0.620 3.020 0.820 ;
        RECT  3.820 0.400 4.020 0.820 ;
        RECT  4.860 0.400 5.060 0.820 ;
        RECT  2.740 0.660 5.060 0.820 ;
        RECT  0.180 1.480 1.500 1.740 ;
        RECT  1.220 1.480 1.500 2.100 ;
        RECT  0.180 1.480 0.460 2.100 ;
        RECT  1.220 1.900 5.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END AOI31M4HM

MACRO AOI31M2HM
    CLASS CORE ;
    FOREIGN AOI31M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.820 1.680 1.290 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.740 1.140 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.340 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.330 1.290 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.753  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.140 1.520 2.700 1.740 ;
        RECT  2.490 0.480 2.700 1.740 ;
        RECT  1.580 0.480 2.700 0.640 ;
        RECT  0.140 1.520 0.420 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.220 -0.140 2.500 0.320 ;
        RECT  0.300 -0.140 0.500 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 1.900 2.020 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI31M2HM

MACRO AOI31M1HM
    CLASS CORE ;
    FOREIGN AOI31M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.820 1.680 1.260 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.740 1.140 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.340 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.330 1.290 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.589  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.140 1.580 2.700 1.740 ;
        RECT  2.490 0.480 2.700 1.740 ;
        RECT  1.580 0.480 2.700 0.640 ;
        RECT  0.140 1.580 0.340 1.970 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.220 -0.140 2.500 0.320 ;
        RECT  0.300 -0.140 0.500 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 1.900 2.060 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI31M1HM

MACRO AOI31M0HM
    CLASS CORE ;
    FOREIGN AOI31M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.820 1.720 1.290 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.740 1.140 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.340 ;
        END
    END A3
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.330 1.290 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.503  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.140 1.580 2.700 1.740 ;
        RECT  2.490 0.480 2.700 1.740 ;
        RECT  1.580 0.480 2.700 0.640 ;
        RECT  0.140 1.580 0.340 2.060 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.220 -0.140 2.500 0.320 ;
        RECT  0.300 -0.140 0.500 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 1.900 2.060 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI31M0HM

MACRO AOI22M8HM
    CLASS CORE ;
    FOREIGN AOI22M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.656  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.080 3.500 1.280 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.420 ;
        LAYER ME1 ;
        RECT  1.160 1.260 3.500 1.420 ;
        RECT  3.300 1.020 3.500 1.420 ;
        RECT  1.160 1.040 1.360 1.420 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.692  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.170 5.500 1.370 ;
        LAYER ME2 ;
        RECT  5.300 1.040 5.500 1.560 ;
        LAYER ME1 ;
        RECT  5.200 1.260 7.760 1.420 ;
        RECT  7.120 1.120 7.760 1.420 ;
        RECT  5.200 1.120 5.840 1.420 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.060 0.800 8.340 1.160 ;
        RECT  4.620 0.800 8.340 0.960 ;
        RECT  6.160 0.800 6.800 1.100 ;
        RECT  4.620 0.800 4.900 1.160 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 1.080 4.240 1.240 ;
        RECT  3.660 0.680 3.820 1.240 ;
        RECT  2.930 0.680 3.820 0.840 ;
        RECT  1.520 0.940 3.090 1.100 ;
        RECT  2.930 0.680 3.090 1.100 ;
        RECT  1.520 0.700 1.680 1.100 ;
        RECT  0.500 0.700 1.680 0.860 ;
        RECT  0.500 0.700 0.700 1.380 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.128  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.740 1.580 8.700 1.740 ;
        RECT  8.500 0.480 8.700 1.740 ;
        RECT  3.980 0.480 8.700 0.640 ;
        RECT  2.590 0.360 4.140 0.520 ;
        RECT  1.830 0.480 2.750 0.640 ;
        RECT  1.100 0.360 1.990 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.260 -0.140 8.540 0.320 ;
        RECT  6.340 -0.140 6.620 0.320 ;
        RECT  4.300 -0.140 4.580 0.320 ;
        RECT  2.150 -0.140 2.430 0.320 ;
        RECT  0.300 -0.140 0.580 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 4.500 1.740 ;
        RECT  4.300 1.580 4.500 2.060 ;
        RECT  0.140 1.580 0.340 1.910 ;
        RECT  4.300 1.900 8.700 2.060 ;
        RECT  8.420 1.900 8.700 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.140 ;
    END
END AOI22M8HM

MACRO AOI22M4HM
    CLASS CORE ;
    FOREIGN AOI22M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.690  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.170 3.500 1.370 ;
        LAYER ME2 ;
        RECT  3.300 1.040 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.120 1.120 3.760 1.420 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.798  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.080 1.500 1.280 ;
        LAYER ME2 ;
        RECT  1.300 0.810 1.500 1.420 ;
        LAYER ME1 ;
        RECT  0.960 1.040 1.580 1.420 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.060 0.800 4.340 1.220 ;
        RECT  2.680 0.800 4.340 0.960 ;
        RECT  2.680 0.800 2.880 1.220 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.740 1.060 2.280 1.260 ;
        RECT  1.740 0.680 1.900 1.260 ;
        RECT  0.500 0.680 1.900 0.840 ;
        RECT  0.500 0.680 0.700 1.380 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.008  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.820 1.580 4.700 1.740 ;
        RECT  4.500 0.480 4.700 1.740 ;
        RECT  2.060 0.480 4.700 0.640 ;
        RECT  1.100 0.360 2.220 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.260 -0.140 4.540 0.320 ;
        RECT  2.380 -0.140 2.660 0.320 ;
        RECT  0.300 -0.140 0.580 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 2.620 1.740 ;
        RECT  2.340 1.580 2.620 2.060 ;
        RECT  0.140 1.580 0.340 1.900 ;
        RECT  2.340 1.900 4.700 2.060 ;
        RECT  4.420 1.900 4.700 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AOI22M4HM

MACRO AOI22M2HM
    CLASS CORE ;
    FOREIGN AOI22M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.600 1.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 0.840 2.300 1.240 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.750 1.100 1.420 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.250 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.602  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.580 2.700 1.740 ;
        RECT  2.500 0.520 2.700 1.740 ;
        RECT  1.660 0.520 2.700 0.680 ;
        RECT  1.660 0.340 1.820 0.680 ;
        RECT  1.080 0.340 1.820 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.060 -0.140 2.340 0.320 ;
        RECT  0.220 -0.140 0.420 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 1.380 1.740 ;
        RECT  1.180 1.580 1.380 2.060 ;
        RECT  0.140 1.580 0.340 2.020 ;
        RECT  1.180 1.900 2.580 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI22M2HM

MACRO AOI22M1HM
    CLASS CORE ;
    FOREIGN AOI22M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.840 1.540 1.370 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 1.980 1.370 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.850 0.840 1.100 1.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.600 1.190 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.372  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.520 1.620 2.300 1.960 ;
        RECT  2.140 0.520 2.300 1.960 ;
        RECT  1.040 0.520 2.300 0.680 ;
        RECT  1.040 0.400 1.410 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  0.540 1.640 0.820 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.180 -0.140 0.380 0.580 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.400 1.050 1.920 2.400 ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.050 ;
        RECT  0.000 0.000 0.400 1.140 ;
        RECT  1.920 0.000 2.400 1.140 ;
    END
END AOI22M1HM

MACRO AOI22M0HM
    CLASS CORE ;
    FOREIGN AOI22M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.280 0.840 1.540 1.370 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 1.980 1.370 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.850 0.840 1.100 1.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.600 1.190 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.303  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.520 1.620 2.300 1.960 ;
        RECT  2.140 0.520 2.300 1.960 ;
        RECT  1.040 0.520 2.300 0.680 ;
        RECT  1.040 0.340 1.410 0.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  0.540 1.640 0.820 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.180 -0.140 0.380 0.560 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI22M0HM

MACRO AOI22B20M8HM
    CLASS CORE ;
    FOREIGN AOI22B20M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.692  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.170 4.700 1.370 ;
        LAYER ME2 ;
        RECT  4.500 1.040 4.700 1.560 ;
        LAYER ME1 ;
        RECT  4.400 1.260 6.960 1.420 ;
        RECT  6.320 1.120 6.960 1.420 ;
        RECT  4.400 1.120 5.040 1.420 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.260 0.800 7.540 1.160 ;
        RECT  3.820 0.800 7.540 0.960 ;
        RECT  5.360 0.800 6.000 1.100 ;
        RECT  3.820 0.800 4.100 1.160 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.820 1.060 1.100 1.560 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.800 0.340 1.300 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.995  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.940 1.580 7.900 1.740 ;
        RECT  7.700 0.480 7.900 1.740 ;
        RECT  1.820 0.480 7.900 0.640 ;
        RECT  2.940 0.360 3.220 0.640 ;
        RECT  1.820 0.340 2.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  2.940 1.900 3.220 2.540 ;
        RECT  1.900 1.820 2.180 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.460 -0.140 7.740 0.320 ;
        RECT  5.540 -0.140 5.820 0.320 ;
        RECT  3.500 -0.140 3.780 0.320 ;
        RECT  2.380 -0.140 2.660 0.320 ;
        RECT  1.300 -0.140 1.580 0.500 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.300 0.860 0.900 ;
        RECT  0.500 0.740 1.520 0.900 ;
        RECT  1.360 0.860 3.300 1.020 ;
        RECT  0.500 0.740 0.660 2.060 ;
        RECT  0.500 1.900 1.280 2.060 ;
        RECT  1.340 1.420 2.660 1.580 ;
        RECT  2.460 1.580 3.700 1.740 ;
        RECT  3.500 1.580 3.700 2.060 ;
        RECT  3.500 1.900 7.900 2.060 ;
        RECT  7.620 1.900 7.900 2.100 ;
        LAYER VTPH ;
        RECT  1.040 1.060 2.960 2.400 ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.060 ;
        RECT  0.000 0.000 1.040 1.140 ;
        RECT  2.960 0.000 8.000 1.140 ;
    END
END AOI22B20M8HM

MACRO AOI22B20M4HM
    CLASS CORE ;
    FOREIGN AOI22B20M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.260 4.240 1.420 ;
        RECT  3.600 1.120 4.240 1.420 ;
        RECT  2.500 0.840 2.700 1.420 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 0.800 4.700 1.320 ;
        RECT  3.100 0.800 4.700 0.960 ;
        RECT  3.100 0.800 3.380 1.100 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.040 1.260 1.320 ;
        RECT  0.900 1.040 1.100 1.600 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.040 0.740 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.907  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 1.580 5.100 1.740 ;
        RECT  4.900 0.480 5.100 1.740 ;
        RECT  2.260 0.480 5.100 0.640 ;
        RECT  2.260 0.330 2.460 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  2.220 1.900 2.500 2.540 ;
        RECT  0.420 1.780 0.620 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.660 -0.140 4.940 0.320 ;
        RECT  2.840 -0.140 3.120 0.320 ;
        RECT  1.700 -0.140 1.980 0.520 ;
        RECT  1.220 -0.140 1.500 0.520 ;
        RECT  0.220 -0.140 0.420 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.760 0.300 0.920 0.840 ;
        RECT  0.760 0.680 1.660 0.840 ;
        RECT  1.500 1.080 2.340 1.280 ;
        RECT  1.500 0.680 1.660 1.670 ;
        RECT  1.280 1.510 1.660 1.670 ;
        RECT  1.280 1.510 1.440 2.100 ;
        RECT  1.860 1.580 2.980 1.740 ;
        RECT  2.780 1.580 2.980 2.060 ;
        RECT  2.780 1.900 5.100 2.060 ;
        RECT  1.860 1.580 2.060 2.080 ;
        RECT  1.700 1.880 2.060 2.080 ;
        RECT  4.820 1.900 5.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END AOI22B20M4HM

MACRO AOI22B20M2HM
    CLASS CORE ;
    FOREIGN AOI22B20M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        ANTENNAGATEAREA 0.059  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 7.252  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.140 1.500 1.340 ;
        LAYER ME2 ;
        RECT  1.300 1.040 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.000 1.080 1.500 1.400 ;
        END
    END NA2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.320 1.400 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.750 3.100 1.360 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.720 1.320 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.501  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 1.580 2.700 1.740 ;
        RECT  2.500 0.340 2.700 1.740 ;
        RECT  1.860 0.340 2.700 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.220 1.900 1.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.880 -0.140 3.100 0.460 ;
        RECT  1.300 -0.140 1.580 0.520 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.410 1.100 0.570 ;
        RECT  0.940 0.410 1.100 0.840 ;
        RECT  0.940 0.680 1.820 0.840 ;
        RECT  1.660 0.680 1.820 1.740 ;
        RECT  0.420 1.580 1.820 1.740 ;
        RECT  0.420 1.580 0.620 2.080 ;
        RECT  1.700 1.900 3.100 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AOI22B20M2HM

MACRO AOI22B20M1HM
    CLASS CORE ;
    FOREIGN AOI22B20M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        ANTENNAGATEAREA 0.059  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.367  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.140 1.100 1.340 ;
        LAYER ME2 ;
        RECT  0.900 1.040 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.900 1.080 1.300 1.400 ;
        END
    END NA2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.050 0.800 2.320 1.250 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.620 3.100 1.400 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.680 1.200 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.442  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.180 1.580 2.700 1.740 ;
        RECT  2.500 0.300 2.700 1.740 ;
        RECT  1.860 0.300 2.700 0.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.100 1.900 1.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.880 -0.140 3.100 0.460 ;
        RECT  1.300 -0.140 1.580 0.520 ;
        RECT  0.140 -0.140 0.340 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.430 1.070 0.590 ;
        RECT  0.910 0.430 1.070 0.840 ;
        RECT  0.910 0.680 1.740 0.840 ;
        RECT  1.580 0.680 1.740 1.740 ;
        RECT  0.300 1.580 1.740 1.740 ;
        RECT  0.300 1.580 0.500 2.070 ;
        RECT  1.620 1.900 3.100 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AOI22B20M1HM

MACRO AOI22B20M0HM
    CLASS CORE ;
    FOREIGN AOI22B20M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        ANTENNAGATEAREA 0.059  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.367  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.140 1.100 1.340 ;
        LAYER ME2 ;
        RECT  0.900 1.040 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.900 1.080 1.300 1.400 ;
        END
    END NA2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.320 1.230 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.800 3.100 1.360 ;
        END
    END B2
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.059  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.680 1.180 ;
        END
    END NA1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.180 1.580 2.700 1.740 ;
        RECT  2.500 0.300 2.700 1.740 ;
        RECT  1.860 0.300 2.700 0.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  1.100 1.900 1.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.880 -0.140 3.100 0.460 ;
        RECT  1.300 -0.140 1.580 0.520 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 0.410 1.030 0.570 ;
        RECT  0.870 0.410 1.030 0.840 ;
        RECT  0.870 0.680 1.740 0.840 ;
        RECT  1.580 0.680 1.740 1.740 ;
        RECT  0.300 1.580 1.740 1.740 ;
        RECT  0.300 1.580 0.500 2.070 ;
        RECT  1.620 1.900 3.100 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AOI22B20M0HM

MACRO AOI222M8HM
    CLASS CORE ;
    FOREIGN AOI222M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  11.840 0.800 12.480 1.100 ;
        RECT  9.760 0.800 12.480 0.960 ;
        RECT  9.760 0.800 10.400 1.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.300 1.260 12.980 1.420 ;
        RECT  12.700 1.080 12.980 1.420 ;
        RECT  10.800 1.120 11.440 1.420 ;
        RECT  9.300 0.840 9.500 1.420 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.680 0.800 8.320 1.100 ;
        RECT  5.600 0.800 8.320 0.960 ;
        RECT  5.600 0.800 6.240 1.100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.100 1.260 8.780 1.420 ;
        RECT  8.500 0.840 8.780 1.420 ;
        RECT  6.640 1.120 7.280 1.420 ;
        RECT  5.100 1.080 5.380 1.420 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.040 0.800 3.680 1.100 ;
        RECT  0.960 0.800 3.680 0.960 ;
        RECT  0.960 0.800 1.600 1.100 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.260 4.180 1.420 ;
        RECT  3.900 1.080 4.180 1.420 ;
        RECT  2.000 1.120 2.640 1.420 ;
        RECT  0.500 0.840 0.700 1.420 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.141  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  9.380 1.580 13.500 1.740 ;
        RECT  13.300 0.480 13.500 1.740 ;
        RECT  1.100 0.480 13.500 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 13.600 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 13.600 0.140 ;
        RECT  12.900 -0.140 13.180 0.320 ;
        RECT  10.980 -0.140 11.260 0.320 ;
        RECT  8.900 -0.140 9.180 0.320 ;
        RECT  6.820 -0.140 7.100 0.320 ;
        RECT  4.900 -0.140 5.180 0.320 ;
        RECT  4.100 -0.140 4.380 0.320 ;
        RECT  2.180 -0.140 2.460 0.320 ;
        RECT  0.340 -0.140 0.540 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.580 1.580 8.700 1.740 ;
        RECT  4.700 1.900 13.380 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 13.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 13.600 1.140 ;
    END
END AOI222M8HM

MACRO AOI222M4HM
    CLASS CORE ;
    FOREIGN AOI222M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.900 1.210 6.240 1.370 ;
        RECT  5.600 1.120 6.240 1.370 ;
        RECT  4.900 1.210 5.100 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.800 6.700 1.180 ;
        RECT  5.100 0.800 6.700 0.960 ;
        RECT  5.100 0.800 5.380 1.040 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.260 4.160 1.420 ;
        RECT  3.520 1.120 4.160 1.420 ;
        RECT  2.500 0.840 2.700 1.420 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.440 0.800 4.700 1.220 ;
        RECT  3.020 0.800 4.700 0.960 ;
        RECT  3.020 0.800 3.300 1.040 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.220 1.600 1.380 ;
        RECT  0.960 1.120 1.600 1.380 ;
        RECT  0.100 0.840 0.300 1.380 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.860 0.800 2.300 1.160 ;
        RECT  0.460 0.800 2.300 0.960 ;
        RECT  0.460 0.800 0.740 1.040 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.069  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.260 1.580 7.100 1.740 ;
        RECT  6.900 0.480 7.100 1.740 ;
        RECT  1.180 0.480 7.100 0.640 ;
        RECT  5.260 1.540 5.540 1.740 ;
        RECT  1.180 0.360 1.380 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.540 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.660 -0.140 6.940 0.320 ;
        RECT  4.740 -0.140 5.020 0.320 ;
        RECT  2.820 -0.140 3.100 0.320 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.340 -0.140 0.540 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.580 4.540 1.740 ;
        RECT  0.660 1.580 0.860 2.060 ;
        RECT  2.620 1.900 7.100 2.060 ;
        RECT  6.820 1.900 7.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END AOI222M4HM

MACRO AOI222M2HM
    CLASS CORE ;
    FOREIGN AOI222M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.450 0.840 0.700 1.250 ;
        END
    END C2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.173  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.140 3.100 1.340 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.900 1.080 3.400 1.400 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.560  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.140 2.300 1.340 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.100 1.080 2.700 1.400 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.800 3.900 1.270 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.750 1.940 1.250 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.960 0.840 1.500 1.160 ;
        END
    END C1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.854  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.140 1.580 4.300 1.740 ;
        RECT  4.100 0.440 4.300 1.740 ;
        RECT  3.300 0.440 4.300 0.600 ;
        RECT  2.140 0.680 3.460 0.840 ;
        RECT  3.300 0.440 3.460 0.840 ;
        RECT  2.140 0.300 2.300 0.840 ;
        RECT  1.140 0.300 2.300 0.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  2.460 0.320 3.140 0.520 ;
        RECT  2.680 -0.140 2.920 0.520 ;
        RECT  0.340 -0.140 0.540 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 2.460 1.740 ;
        RECT  0.140 1.580 0.340 1.900 ;
        RECT  1.580 1.900 4.020 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AOI222M2HM

MACRO AOI222M1HM
    CLASS CORE ;
    FOREIGN AOI222M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.450 0.840 0.700 1.280 ;
        END
    END C2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        ANTENNAGATEAREA 0.095  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.046  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.140 3.100 1.340 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.900 1.080 3.500 1.400 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        ANTENNAGATEAREA 0.095  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.046  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.140 2.300 1.340 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.100 1.080 2.700 1.400 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.800 3.920 1.320 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.760 1.940 1.400 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.960 0.840 1.500 1.200 ;
        END
    END C1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.682  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.580 4.300 1.740 ;
        RECT  4.100 0.340 4.300 1.740 ;
        RECT  3.300 0.340 4.300 0.500 ;
        RECT  2.140 0.680 3.460 0.840 ;
        RECT  3.300 0.340 3.460 0.840 ;
        RECT  2.140 0.300 2.300 0.840 ;
        RECT  1.140 0.300 2.300 0.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  2.460 0.320 3.140 0.520 ;
        RECT  2.680 -0.140 2.920 0.520 ;
        RECT  0.340 -0.140 0.540 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 2.500 1.740 ;
        RECT  0.140 1.580 0.340 1.960 ;
        RECT  1.180 1.580 1.380 1.960 ;
        RECT  1.580 1.900 4.180 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AOI222M1HM

MACRO AOI222M0HM
    CLASS CORE ;
    FOREIGN AOI222M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.328  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.140 2.300 1.340 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.100 1.080 2.700 1.400 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.328  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.140 3.100 1.340 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.900 1.080 3.500 1.400 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 0.840 3.920 1.320 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.800 1.940 1.400 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.000 0.840 1.500 1.200 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.750 1.240 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.614  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.580 4.300 1.740 ;
        RECT  4.100 0.300 4.300 1.740 ;
        RECT  3.300 0.300 4.300 0.460 ;
        RECT  2.140 0.680 3.460 0.840 ;
        RECT  3.300 0.300 3.460 0.840 ;
        RECT  2.140 0.300 2.300 0.840 ;
        RECT  1.140 0.300 2.300 0.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  2.500 0.320 3.140 0.520 ;
        RECT  2.680 -0.140 2.920 0.520 ;
        RECT  0.280 -0.140 0.480 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.580 2.500 1.740 ;
        RECT  0.100 1.580 0.380 1.960 ;
        RECT  1.140 1.580 1.420 1.960 ;
        RECT  1.580 1.900 4.180 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AOI222M0HM

MACRO AOI221M8HM
    CLASS CORE ;
    FOREIGN AOI221M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.000 0.800 10.640 1.100 ;
        RECT  7.920 0.800 10.640 0.960 ;
        RECT  7.920 0.800 8.560 1.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.420 1.260 11.140 1.420 ;
        RECT  10.860 0.840 11.140 1.420 ;
        RECT  8.960 1.120 9.600 1.420 ;
        RECT  7.420 1.060 7.700 1.420 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.360 0.800 6.000 1.100 ;
        RECT  3.280 0.800 6.000 0.960 ;
        RECT  3.280 0.800 3.920 1.100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.536  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.800 1.260 6.440 1.420 ;
        RECT  6.240 1.000 6.440 1.420 ;
        RECT  4.320 1.120 4.960 1.420 ;
        RECT  2.800 0.840 3.100 1.420 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.476  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.780 0.840 2.260 1.240 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.092  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.540 1.580 11.500 1.740 ;
        RECT  11.300 0.480 11.500 1.740 ;
        RECT  0.740 0.480 11.500 0.640 ;
        RECT  10.180 0.390 10.460 0.640 ;
        RECT  8.100 0.390 8.380 0.640 ;
        RECT  5.540 0.390 5.820 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.600 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.600 0.140 ;
        RECT  11.060 -0.140 11.340 0.320 ;
        RECT  9.140 -0.140 9.420 0.320 ;
        RECT  7.220 -0.140 7.500 0.320 ;
        RECT  6.420 -0.140 6.700 0.320 ;
        RECT  4.500 -0.140 4.780 0.320 ;
        RECT  2.520 -0.140 2.800 0.320 ;
        RECT  1.340 -0.140 1.620 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.340 1.580 6.900 1.740 ;
        RECT  0.340 1.580 0.560 2.100 ;
        RECT  1.420 1.580 1.620 2.100 ;
        RECT  2.460 1.580 2.660 2.100 ;
        RECT  2.900 1.900 11.500 2.060 ;
        RECT  11.220 1.900 11.500 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 11.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.600 1.140 ;
    END
END AOI221M8HM

MACRO AOI221M4HM
    CLASS CORE ;
    FOREIGN AOI221M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.210 5.440 1.370 ;
        RECT  4.800 1.120 5.440 1.370 ;
        RECT  4.100 1.210 4.300 1.560 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.700 0.800 5.900 1.320 ;
        RECT  4.300 0.800 5.900 0.960 ;
        RECT  4.300 0.800 4.580 1.040 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.240 1.210 3.900 1.370 ;
        RECT  3.700 0.840 3.900 1.370 ;
        RECT  2.240 1.120 2.880 1.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.100 0.800 3.380 1.040 ;
        RECT  1.700 0.800 3.380 0.960 ;
        RECT  1.700 0.800 1.980 1.320 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.239  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 0.900 1.270 1.320 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.021  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.460 1.580 6.300 1.740 ;
        RECT  6.100 0.480 6.300 1.740 ;
        RECT  0.900 0.480 6.300 0.640 ;
        RECT  5.020 0.360 5.220 0.640 ;
        RECT  4.460 1.540 4.740 1.740 ;
        RECT  2.460 0.360 2.660 0.640 ;
        RECT  0.900 0.300 1.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  0.860 1.900 1.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.860 -0.140 6.140 0.320 ;
        RECT  4.100 -0.140 4.380 0.320 ;
        RECT  3.300 -0.140 3.580 0.320 ;
        RECT  1.480 -0.140 1.760 0.320 ;
        RECT  0.380 -0.140 0.580 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.300 1.580 3.780 1.740 ;
        RECT  1.860 1.900 6.300 2.060 ;
        RECT  6.020 1.900 6.300 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
    END
END AOI221M4HM

MACRO AOI221M2HM
    CLASS CORE ;
    FOREIGN AOI221M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.173  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.140 2.700 1.340 ;
        LAYER ME2 ;
        RECT  2.500 1.040 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.200 1.080 2.700 1.400 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.708  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.160 1.100 1.360 ;
        LAYER ME2 ;
        RECT  0.900 1.040 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.860 1.000 1.140 1.420 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.560  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.080 1.900 1.400 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.750 3.100 1.360 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.040 0.440 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.600  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.620 1.580 3.500 1.740 ;
        RECT  3.300 0.300 3.500 1.740 ;
        RECT  2.580 0.300 3.500 0.460 ;
        RECT  0.680 0.680 2.740 0.840 ;
        RECT  2.580 0.300 2.740 0.840 ;
        RECT  0.680 0.370 0.840 0.840 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.140 -0.140 2.420 0.520 ;
        RECT  1.460 -0.140 1.740 0.520 ;
        RECT  0.140 -0.140 0.340 0.690 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.580 1.900 1.980 2.060 ;
        RECT  1.100 1.580 2.380 1.740 ;
        RECT  2.180 1.580 2.380 2.060 ;
        RECT  2.180 1.900 3.500 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI221M2HM

MACRO AOI221M1HM
    CLASS CORE ;
    FOREIGN AOI221M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.084  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.200 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.860 0.800 3.100 1.250 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.380 0.840 2.700 1.200 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.100 1.200 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.095  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.600 1.200 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.520  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.600 1.580 3.500 1.740 ;
        RECT  3.300 0.300 3.500 1.740 ;
        RECT  2.580 0.300 3.500 0.460 ;
        RECT  0.700 0.480 2.740 0.640 ;
        RECT  2.580 0.300 2.740 0.640 ;
        RECT  0.700 0.340 0.980 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  0.100 1.700 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  1.580 -0.140 2.380 0.320 ;
        RECT  0.140 -0.140 0.340 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.740 1.420 2.020 1.660 ;
        RECT  0.580 1.500 2.020 1.660 ;
        RECT  1.140 1.900 3.480 2.060 ;
        RECT  3.200 1.900 3.480 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.060 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.060 ;
    END
END AOI221M1HM

MACRO AOI221M0HM
    CLASS CORE ;
    FOREIGN AOI221M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.560 1.180 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.620 3.100 1.420 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.380 0.840 2.700 1.200 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.100 1.200 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.620 1.200 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.486  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.600 1.580 3.500 1.740 ;
        RECT  3.300 0.300 3.500 1.740 ;
        RECT  2.580 0.300 3.500 0.460 ;
        RECT  0.700 0.480 2.740 0.640 ;
        RECT  2.580 0.300 2.740 0.640 ;
        RECT  0.700 0.370 0.980 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  0.100 1.600 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  1.620 -0.140 2.380 0.320 ;
        RECT  0.140 -0.140 0.340 0.470 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.740 1.420 2.020 1.660 ;
        RECT  0.580 1.500 2.020 1.660 ;
        RECT  1.140 1.900 3.480 2.060 ;
        RECT  3.200 1.900 3.480 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.060 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.060 ;
    END
END AOI221M0HM

MACRO AOI21M8HM
    CLASS CORE ;
    FOREIGN AOI21M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        ANTENNAGATEAREA 0.580  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.727  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.300 1.170 5.500 1.370 ;
        LAYER ME2 ;
        RECT  5.300 1.040 5.500 1.560 ;
        LAYER ME1 ;
        RECT  3.180 1.260 5.780 1.420 ;
        RECT  5.140 1.120 5.780 1.420 ;
        RECT  3.180 1.120 3.820 1.420 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.580  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.140 0.800 6.300 1.260 ;
        RECT  2.500 0.800 6.300 0.960 ;
        RECT  4.160 0.800 4.800 1.100 ;
        RECT  2.500 0.800 2.820 1.220 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.620 0.900 1.300 1.230 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.109  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.580 6.700 1.740 ;
        RECT  6.500 0.480 6.700 1.740 ;
        RECT  0.580 0.480 6.700 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  1.740 1.900 2.020 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.300 -0.140 6.580 0.320 ;
        RECT  4.340 -0.140 4.620 0.320 ;
        RECT  2.340 -0.140 2.620 0.320 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 1.580 2.540 1.740 ;
        RECT  2.260 1.580 2.540 2.060 ;
        RECT  2.260 1.900 6.700 2.060 ;
        RECT  0.220 1.580 0.420 2.100 ;
        RECT  1.260 1.580 1.460 2.100 ;
        RECT  6.420 1.900 6.700 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
    END
END AOI21M8HM

MACRO AOI21M6HM
    CLASS CORE ;
    FOREIGN AOI21M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.433  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.500 0.800 4.700 1.250 ;
        RECT  2.520 0.800 4.700 0.960 ;
        RECT  2.520 0.800 2.800 1.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.433  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 1.260 4.240 1.420 ;
        RECT  3.440 1.120 4.240 1.420 ;
        RECT  2.100 0.840 2.300 1.420 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.379  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.810 1.300 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.493  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.180 1.580 5.100 1.740 ;
        RECT  4.900 0.480 5.100 1.740 ;
        RECT  1.140 0.480 5.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.180 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  3.700 -0.140 3.980 0.320 ;
        RECT  1.740 -0.140 2.020 0.320 ;
        RECT  0.700 -0.140 0.900 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 1.580 1.940 1.740 ;
        RECT  1.740 1.580 1.940 2.060 ;
        RECT  1.740 1.900 5.100 2.060 ;
        RECT  4.820 1.900 5.100 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END AOI21M6HM

MACRO AOI21M4HM
    CLASS CORE ;
    FOREIGN AOI21M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.260 2.640 1.420 ;
        RECT  2.000 1.120 2.640 1.420 ;
        RECT  0.900 0.840 1.100 1.420 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.800 3.100 1.210 ;
        RECT  1.480 0.800 3.100 0.960 ;
        RECT  1.480 0.800 1.760 1.100 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.660 1.160 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.907  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 1.580 3.500 1.740 ;
        RECT  3.300 0.480 3.500 1.740 ;
        RECT  0.660 0.480 3.500 0.640 ;
        RECT  0.660 0.330 0.860 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  1.240 -0.140 1.520 0.320 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 1.380 1.740 ;
        RECT  1.180 1.580 1.380 2.060 ;
        RECT  0.140 1.580 0.340 1.960 ;
        RECT  1.180 1.900 3.500 2.060 ;
        RECT  3.220 1.900 3.500 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI21M4HM

MACRO AOI21M3HM
    CLASS CORE ;
    FOREIGN AOI21M3HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.180 2.640 1.340 ;
        RECT  2.000 1.120 2.640 1.340 ;
        RECT  0.900 0.840 1.100 1.340 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.220  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 0.800 3.100 1.160 ;
        RECT  1.480 0.800 3.100 0.960 ;
        RECT  1.480 0.800 1.760 1.020 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.660 1.200 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.686  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.500 3.500 1.660 ;
        RECT  3.300 0.480 3.500 1.660 ;
        RECT  0.660 0.480 3.500 0.640 ;
        RECT  2.700 1.500 2.980 1.750 ;
        RECT  1.660 1.500 1.940 1.750 ;
        RECT  0.660 0.330 0.860 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.060 -0.140 3.340 0.320 ;
        RECT  1.240 -0.140 1.520 0.320 ;
        RECT  0.140 -0.140 0.340 0.610 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.580 1.380 1.740 ;
        RECT  1.180 1.580 1.380 2.100 ;
        RECT  2.180 1.820 2.460 2.100 ;
        RECT  0.140 1.580 0.340 1.960 ;
        RECT  3.220 1.820 3.500 2.100 ;
        RECT  1.180 1.940 3.500 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI21M3HM

MACRO AOI21M2HM
    CLASS CORE ;
    FOREIGN AOI21M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.180 1.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.320 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 0.840 1.900 1.320 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.671  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.580 2.300 1.740 ;
        RECT  2.100 0.480 2.300 1.740 ;
        RECT  1.400 0.480 2.300 0.640 ;
        RECT  1.400 0.360 1.600 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.960 2.080 2.240 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.960 -0.140 2.240 0.320 ;
        RECT  0.200 -0.140 0.400 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.120 1.900 1.680 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI21M2HM

MACRO AOI21M1HM
    CLASS CORE ;
    FOREIGN AOI21M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.220 1.230 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.420 0.840 0.700 1.320 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 0.840 1.900 1.320 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.505  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.580 2.300 1.740 ;
        RECT  2.100 0.480 2.300 1.740 ;
        RECT  1.400 0.480 2.300 0.640 ;
        RECT  1.400 0.360 1.600 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.960 2.080 2.240 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.960 -0.140 2.240 0.320 ;
        RECT  0.200 -0.140 0.400 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.120 1.900 1.680 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI21M1HM

MACRO AOI21M0HM
    CLASS CORE ;
    FOREIGN AOI21M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.180 1.230 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.350 0.840 0.700 1.280 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.480 1.080 1.900 1.400 ;
        RECT  1.700 0.840 1.900 1.400 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.433  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.720 1.580 2.300 1.740 ;
        RECT  2.100 0.480 2.300 1.740 ;
        RECT  1.400 0.480 2.300 0.640 ;
        RECT  1.400 0.320 1.600 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  1.960 2.080 2.240 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.960 -0.140 2.240 0.320 ;
        RECT  0.200 -0.140 0.400 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.120 1.900 1.680 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI21M0HM

MACRO AOI21B20M8HM
    CLASS CORE ;
    FOREIGN AOI21B20M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.504  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.040 0.800 4.680 1.100 ;
        RECT  2.040 0.800 4.680 0.960 ;
        RECT  2.040 0.800 2.720 1.100 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.200 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.000 1.100 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.190  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.180 1.760 5.500 1.920 ;
        RECT  5.300 0.480 5.500 1.920 ;
        RECT  1.900 0.480 5.500 0.640 ;
        RECT  1.620 0.340 2.060 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.100 2.080 5.380 2.540 ;
        RECT  3.340 2.080 3.620 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  4.460 -0.140 4.740 0.320 ;
        RECT  3.340 -0.140 3.620 0.320 ;
        RECT  2.220 -0.140 2.500 0.320 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.340 0.980 0.540 ;
        RECT  0.780 0.340 0.980 0.820 ;
        RECT  0.780 0.660 1.720 0.820 ;
        RECT  3.160 1.120 3.800 1.420 ;
        RECT  4.940 0.980 5.100 1.420 ;
        RECT  1.560 1.260 5.100 1.420 ;
        RECT  1.560 0.660 1.720 1.920 ;
        RECT  0.100 1.720 1.720 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END AOI21B20M8HM

MACRO AOI21B20M4HM
    CLASS CORE ;
    FOREIGN AOI21B20M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.568  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.140 1.760 3.500 1.920 ;
        RECT  3.300 0.680 3.500 1.920 ;
        RECT  1.860 0.680 3.500 0.840 ;
        RECT  2.740 0.330 2.940 0.840 ;
        RECT  1.860 0.380 2.020 0.840 ;
        RECT  1.620 0.380 2.020 0.540 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        ANTENNAGATEAREA 0.252  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.837  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.030 2.300 1.230 ;
        LAYER ME2 ;
        RECT  2.100 0.840 2.300 1.360 ;
        LAYER ME1 ;
        RECT  2.000 1.030 2.640 1.280 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.080 0.600 1.560 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.840 1.040 1.160 1.500 ;
        END
    END NA2
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.520 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        RECT  1.140 -0.140 1.420 0.540 ;
        RECT  0.140 -0.140 0.340 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.060 2.080 3.340 2.540 ;
        RECT  1.140 2.080 1.420 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.660 0.330 0.860 0.860 ;
        RECT  0.660 0.700 1.700 0.860 ;
        RECT  2.920 1.020 3.080 1.600 ;
        RECT  1.540 1.440 3.080 1.600 ;
        RECT  1.540 0.700 1.700 1.920 ;
        RECT  0.100 1.720 1.700 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AOI21B20M4HM

MACRO AOI21B20M2HM
    CLASS CORE ;
    FOREIGN AOI21B20M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.050 0.990 2.300 1.560 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.510 1.200 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.040 1.150 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.379  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.720 2.700 2.060 ;
        RECT  2.500 0.620 2.700 2.060 ;
        RECT  1.980 0.620 2.700 0.820 ;
        RECT  1.980 0.320 2.180 0.820 ;
        RECT  1.740 0.320 2.180 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.940 2.080 1.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.340 -0.140 2.540 0.460 ;
        RECT  1.180 -0.140 1.460 0.520 ;
        RECT  0.100 -0.140 0.380 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.300 0.900 0.840 ;
        RECT  0.680 0.680 1.820 0.840 ;
        RECT  1.660 0.680 1.820 1.920 ;
        RECT  0.100 1.720 1.820 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B20M2HM

MACRO AOI21B20M1HM
    CLASS CORE ;
    FOREIGN AOI21B20M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.050 1.040 2.320 1.560 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.040 1.100 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.294  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.790 2.700 1.990 ;
        RECT  2.500 0.620 2.700 1.990 ;
        RECT  1.980 0.620 2.700 0.820 ;
        RECT  1.980 0.300 2.180 0.820 ;
        RECT  1.780 0.300 2.180 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.940 2.080 1.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.420 -0.140 2.620 0.460 ;
        RECT  1.180 -0.140 1.460 0.520 ;
        RECT  0.140 -0.140 0.340 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.340 1.000 0.540 ;
        RECT  0.800 0.340 1.000 0.840 ;
        RECT  0.800 0.680 1.820 0.840 ;
        RECT  1.660 0.680 1.820 1.920 ;
        RECT  0.100 1.720 1.820 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B20M1HM

MACRO AOI21B20M0HM
    CLASS CORE ;
    FOREIGN AOI21B20M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.050 1.040 2.320 1.560 ;
        END
    END B
    PIN NA1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.250 ;
        END
    END NA1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.040 1.150 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.250  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.790 2.700 1.990 ;
        RECT  2.500 0.620 2.700 1.990 ;
        RECT  1.980 0.620 2.700 0.820 ;
        RECT  1.980 0.300 2.180 0.820 ;
        RECT  1.780 0.300 2.180 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.940 2.080 1.700 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.420 -0.140 2.620 0.460 ;
        RECT  1.180 -0.140 1.460 0.520 ;
        RECT  0.100 -0.140 0.380 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.340 0.990 0.540 ;
        RECT  0.790 0.340 0.990 0.840 ;
        RECT  0.790 0.680 1.820 0.840 ;
        RECT  1.660 0.680 1.820 1.920 ;
        RECT  0.100 1.720 1.820 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B20M0HM

MACRO AOI21B10M8HM
    CLASS CORE ;
    FOREIGN AOI21B10M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.553  LAYER ME2  ;
        ANTENNAGATEAREA 0.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.970  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.120 6.300 1.320 ;
        LAYER ME2 ;
        RECT  6.100 1.040 6.300 1.560 ;
        LAYER ME1 ;
        RECT  3.720 1.260 6.440 1.420 ;
        RECT  5.800 1.120 6.440 1.420 ;
        RECT  3.720 1.120 4.360 1.420 ;
        END
    END A1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.935  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.040 0.700 1.380 ;
        END
    END NA2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.485  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.870 2.660 1.070 ;
        RECT  1.180 0.870 1.560 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.753  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.340 1.580 7.500 1.740 ;
        RECT  7.300 0.480 7.500 1.740 ;
        RECT  1.260 0.480 7.500 0.640 ;
        RECT  3.900 0.330 4.180 0.640 ;
        RECT  2.380 0.310 2.580 0.640 ;
        RECT  1.260 0.310 1.460 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  2.300 2.080 2.580 2.540 ;
        RECT  1.260 1.780 1.460 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.860 -0.140 7.140 0.320 ;
        RECT  4.940 -0.140 5.220 0.320 ;
        RECT  2.960 -0.140 3.240 0.320 ;
        RECT  1.780 -0.140 2.060 0.320 ;
        RECT  0.660 -0.140 0.940 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.370 0.320 0.820 ;
        RECT  0.160 0.660 1.020 0.820 ;
        RECT  3.280 0.800 6.880 0.960 ;
        RECT  4.600 0.800 5.480 1.100 ;
        RECT  6.720 0.800 6.880 1.320 ;
        RECT  3.280 0.800 3.440 1.360 ;
        RECT  3.020 1.130 3.440 1.360 ;
        RECT  0.860 1.440 3.180 1.600 ;
        RECT  3.020 1.130 3.180 1.600 ;
        RECT  0.860 0.660 1.020 1.740 ;
        RECT  0.160 1.580 1.020 1.740 ;
        RECT  0.160 1.580 0.320 2.060 ;
        RECT  1.700 1.760 3.140 1.920 ;
        RECT  2.860 1.900 7.340 2.060 ;
        LAYER VTPH ;
        RECT  1.060 0.910 3.300 2.400 ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 0.910 ;
        RECT  0.000 0.000 1.060 1.140 ;
        RECT  3.300 0.000 7.600 1.140 ;
    END
END AOI21B10M8HM

MACRO AOI21B10M4HM
    CLASS CORE ;
    FOREIGN AOI21B10M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.290  LAYER ME1  ;
        ANTENNAGATEAREA 0.290  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.737  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.120 3.500 1.320 ;
        LAYER ME2 ;
        RECT  3.300 1.040 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.960 1.120 3.680 1.370 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.252  LAYER ME1  ;
        ANTENNAGATEAREA 0.252  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.837  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.120 1.500 1.320 ;
        LAYER ME2 ;
        RECT  1.300 1.040 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.180 1.120 1.820 1.370 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.904  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.540 4.700 1.720 ;
        RECT  4.500 0.480 4.700 1.720 ;
        RECT  1.180 0.480 4.700 0.640 ;
        RECT  3.700 1.540 3.980 1.780 ;
        RECT  2.660 1.540 2.940 1.780 ;
        RECT  1.180 0.310 1.380 0.640 ;
        END
    END Z
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.040 0.700 1.380 ;
        END
    END NA2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.060 -0.140 4.340 0.320 ;
        RECT  2.300 -0.140 2.580 0.320 ;
        RECT  1.700 -0.140 1.980 0.320 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.160 0.300 0.320 0.820 ;
        RECT  0.160 0.660 1.020 0.820 ;
        RECT  0.860 0.800 4.080 0.960 ;
        RECT  2.500 0.800 2.780 1.280 ;
        RECT  3.920 0.800 4.080 1.320 ;
        RECT  0.860 0.660 1.020 1.740 ;
        RECT  0.160 1.580 1.020 1.740 ;
        RECT  0.160 1.580 0.320 2.060 ;
        RECT  1.180 1.540 2.420 1.740 ;
        RECT  1.180 1.540 1.380 1.900 ;
        RECT  2.100 1.540 2.420 2.100 ;
        RECT  3.180 1.900 3.460 2.100 ;
        RECT  4.220 1.900 4.500 2.100 ;
        RECT  2.100 1.940 4.500 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AOI21B10M4HM

MACRO AOI21B10M2HM
    CLASS CORE ;
    FOREIGN AOI21B10M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.259  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.120 1.960 1.370 ;
        END
    END A1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.899  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.120 0.300 1.320 ;
        LAYER ME2 ;
        RECT  0.100 1.040 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.080 0.980 0.420 1.420 ;
        END
    END NA2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.126  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.140 1.610 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.574  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 1.540 2.700 1.740 ;
        RECT  2.500 0.480 2.700 1.740 ;
        RECT  1.980 0.480 2.700 0.640 ;
        RECT  1.200 0.340 2.140 0.500 ;
        RECT  1.620 1.540 1.920 1.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.300 -0.140 2.580 0.320 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.320 0.380 0.820 ;
        RECT  0.100 0.660 1.820 0.820 ;
        RECT  1.600 0.800 2.280 0.960 ;
        RECT  2.120 0.800 2.280 1.320 ;
        RECT  0.580 0.660 0.740 1.740 ;
        RECT  0.100 1.580 0.740 1.740 ;
        RECT  0.100 1.580 0.380 2.080 ;
        RECT  1.100 1.840 1.420 2.080 ;
        RECT  2.140 1.900 2.500 2.080 ;
        RECT  1.100 1.920 2.500 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B10M2HM

MACRO AOI21B10M1HM
    CLASS CORE ;
    FOREIGN AOI21B10M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.899  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.120 0.300 1.320 ;
        LAYER ME2 ;
        RECT  0.100 1.040 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.080 0.980 0.420 1.420 ;
        END
    END NA2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        ANTENNAGATEAREA 0.102  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.639  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.120 1.960 1.370 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.089  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.980 1.140 1.610 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.471  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.540 2.700 1.740 ;
        RECT  2.500 0.480 2.700 1.740 ;
        RECT  2.060 0.480 2.700 0.640 ;
        RECT  1.200 0.340 2.220 0.500 ;
        RECT  1.660 1.540 1.960 1.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.380 -0.140 2.660 0.320 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.320 0.380 0.820 ;
        RECT  0.100 0.660 1.820 0.820 ;
        RECT  1.600 0.800 2.340 0.960 ;
        RECT  2.180 0.800 2.340 1.320 ;
        RECT  0.580 0.660 0.740 1.740 ;
        RECT  0.100 1.580 0.740 1.740 ;
        RECT  0.100 1.580 0.380 2.080 ;
        RECT  1.100 1.840 1.420 2.080 ;
        RECT  2.220 1.900 2.580 2.080 ;
        RECT  1.100 1.920 2.580 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B10M1HM

MACRO AOI21B10M0HM
    CLASS CORE ;
    FOREIGN AOI21B10M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.773  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.100 1.120 0.300 1.320 ;
        LAYER ME2 ;
        RECT  0.100 1.040 0.300 1.560 ;
        LAYER ME1 ;
        RECT  0.080 1.000 0.420 1.420 ;
        END
    END NA2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        ANTENNAGATEAREA 0.080  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.821  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.160 1.900 1.360 ;
        LAYER ME2 ;
        RECT  1.700 1.040 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.140 1.960 1.380 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.000 1.140 1.610 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.405  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 1.580 2.700 1.740 ;
        RECT  2.520 0.500 2.700 1.740 ;
        RECT  2.500 1.240 2.700 1.740 ;
        RECT  2.060 0.500 2.700 0.660 ;
        RECT  1.200 0.360 2.220 0.520 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.380 -0.140 2.660 0.340 ;
        RECT  0.620 -0.140 0.900 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 0.380 0.840 ;
        RECT  0.100 0.680 1.820 0.840 ;
        RECT  1.600 0.820 2.360 0.980 ;
        RECT  2.160 0.820 2.360 1.140 ;
        RECT  0.580 0.680 0.740 1.740 ;
        RECT  0.100 1.580 0.740 1.740 ;
        RECT  0.100 1.580 0.380 2.080 ;
        RECT  1.100 1.900 2.580 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B10M0HM

MACRO AOI21B01M8HM
    CLASS CORE ;
    FOREIGN AOI21B01M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.553  LAYER ME2  ;
        ANTENNAGATEAREA 0.553  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.801  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.100 1.120 6.300 1.320 ;
        LAYER ME2 ;
        RECT  6.100 1.040 6.300 1.560 ;
        LAYER ME1 ;
        RECT  3.820 1.260 6.360 1.420 ;
        RECT  5.720 1.120 6.360 1.420 ;
        RECT  3.820 1.120 4.100 1.420 ;
        END
    END A1
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.935  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.040 0.700 1.380 ;
        END
    END NB
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.553  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.640 0.800 6.800 1.320 ;
        RECT  3.220 0.800 6.800 0.960 ;
        RECT  4.520 0.800 5.480 1.100 ;
        RECT  3.220 0.800 3.500 1.360 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.753  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.580 7.500 1.740 ;
        RECT  7.300 0.480 7.500 1.740 ;
        RECT  1.380 0.480 7.500 0.640 ;
        RECT  3.860 0.330 4.060 0.640 ;
        RECT  2.300 0.310 2.500 0.640 ;
        RECT  1.100 0.340 1.540 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  2.260 1.880 2.540 2.540 ;
        RECT  1.260 1.430 1.460 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  6.780 -0.140 7.060 0.320 ;
        RECT  4.860 -0.140 5.140 0.320 ;
        RECT  2.880 -0.140 3.160 0.320 ;
        RECT  1.700 -0.140 1.980 0.320 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.410 0.340 0.840 ;
        RECT  0.140 0.660 1.060 0.840 ;
        RECT  0.860 0.850 2.580 1.050 ;
        RECT  0.860 0.660 1.060 1.740 ;
        RECT  0.100 1.540 1.060 1.740 ;
        RECT  0.100 1.540 0.380 2.100 ;
        RECT  1.740 1.500 3.060 1.720 ;
        RECT  2.780 1.500 3.060 2.100 ;
        RECT  1.740 1.500 2.020 2.100 ;
        RECT  2.780 1.900 7.220 2.100 ;
        LAYER VTPH ;
        RECT  1.060 0.910 3.220 2.400 ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 0.910 ;
        RECT  0.000 0.000 1.060 1.140 ;
        RECT  3.220 0.000 7.600 1.140 ;
    END
END AOI21B01M8HM

MACRO AOI21B01M4HM
    CLASS CORE ;
    FOREIGN AOI21B01M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.290  LAYER ME1  ;
        ANTENNAGATEAREA 0.290  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.594  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.120 3.500 1.320 ;
        LAYER ME2 ;
        RECT  3.300 1.040 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.000 1.120 3.640 1.370 ;
        END
    END A1
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        ANTENNAGATEAREA 0.101  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.333  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.040 0.700 1.380 ;
        END
    END NB
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.290  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 0.800 4.100 1.320 ;
        RECT  2.500 0.800 4.100 0.960 ;
        RECT  2.500 0.800 2.700 1.360 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.904  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.620 1.540 4.700 1.700 ;
        RECT  4.500 0.480 4.700 1.700 ;
        RECT  1.660 0.480 4.700 0.640 ;
        RECT  1.660 0.330 1.860 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  1.620 1.900 1.900 2.540 ;
        RECT  0.140 1.540 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.060 -0.140 4.340 0.320 ;
        RECT  2.240 -0.140 2.520 0.320 ;
        RECT  1.100 -0.140 1.380 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.310 0.340 0.840 ;
        RECT  0.140 0.660 1.100 0.840 ;
        RECT  0.900 0.960 2.080 1.160 ;
        RECT  0.900 0.660 1.100 1.740 ;
        RECT  0.620 1.540 1.100 1.740 ;
        RECT  1.260 1.540 2.420 1.740 ;
        RECT  2.100 1.540 2.420 2.060 ;
        RECT  2.100 1.900 4.540 2.060 ;
        RECT  1.260 1.540 1.460 2.080 ;
        RECT  1.060 1.900 1.460 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AOI21B01M4HM

MACRO AOI21B01M2HM
    CLASS CORE ;
    FOREIGN AOI21B01M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.275  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.200 1.040 0.700 1.380 ;
        END
    END NB
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.800 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.340 1.400 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.510  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 1.560 2.700 1.720 ;
        RECT  2.500 0.480 2.700 1.720 ;
        RECT  1.340 0.480 2.700 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.780 1.900 1.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.260 -0.140 2.540 0.320 ;
        RECT  0.780 -0.140 1.060 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.300 0.300 0.500 0.860 ;
        RECT  0.300 0.660 1.140 0.860 ;
        RECT  0.940 0.660 1.140 1.740 ;
        RECT  0.300 1.540 1.140 1.740 ;
        RECT  0.300 1.540 0.500 2.060 ;
        RECT  1.300 1.540 1.580 2.100 ;
        RECT  2.340 1.900 2.620 2.100 ;
        RECT  1.300 1.940 2.620 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B01M2HM

MACRO AOI21B01M1HM
    CLASS CORE ;
    FOREIGN AOI21B01M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.778  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.120 0.700 1.320 ;
        LAYER ME2 ;
        RECT  0.500 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.120 1.040 0.700 1.380 ;
        END
    END NB
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.840 1.720 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.340 1.280 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.419  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 1.560 2.700 1.740 ;
        RECT  2.500 0.480 2.700 1.740 ;
        RECT  1.780 0.480 2.700 0.640 ;
        RECT  1.780 1.560 2.070 1.780 ;
        RECT  1.300 0.330 1.950 0.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.260 -0.140 2.540 0.320 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 0.300 0.420 0.860 ;
        RECT  0.220 0.660 1.060 0.860 ;
        RECT  0.860 0.660 1.060 1.740 ;
        RECT  0.220 1.540 1.060 1.740 ;
        RECT  0.220 1.540 0.420 2.060 ;
        RECT  1.260 1.790 1.460 2.100 ;
        RECT  2.340 1.900 2.620 2.100 ;
        RECT  1.260 1.940 2.620 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B01M1HM

MACRO AOI21B01M0HM
    CLASS CORE ;
    FOREIGN AOI21B01M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN NB
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.275  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.420 1.120 0.620 1.320 ;
        LAYER ME2 ;
        RECT  0.420 1.040 0.700 1.560 ;
        LAYER ME1 ;
        RECT  0.120 1.040 0.620 1.380 ;
        END
    END NB
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.220 0.840 1.720 1.200 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.340 1.400 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.364  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.780 1.560 2.700 1.740 ;
        RECT  2.500 0.480 2.700 1.740 ;
        RECT  1.480 0.480 2.700 0.640 ;
        RECT  1.780 1.560 2.060 1.780 ;
        RECT  1.300 0.330 1.640 0.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  0.700 1.900 0.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.260 -0.140 2.540 0.320 ;
        RECT  0.700 -0.140 0.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 0.310 0.420 0.860 ;
        RECT  0.220 0.660 1.060 0.860 ;
        RECT  0.860 0.660 1.060 1.740 ;
        RECT  0.220 1.540 1.060 1.740 ;
        RECT  0.220 1.540 0.420 2.060 ;
        RECT  1.260 1.810 1.460 2.100 ;
        RECT  2.340 1.900 2.620 2.100 ;
        RECT  1.260 1.940 2.620 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AOI21B01M0HM

MACRO AOI211M8HM
    CLASS CORE ;
    FOREIGN AOI211M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.538  LAYER ME1  ;
        ANTENNAGATEAREA 0.538  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.095  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  6.500 1.150 6.700 1.350 ;
        LAYER ME2 ;
        RECT  6.500 1.070 6.700 1.590 ;
        LAYER ME1 ;
        RECT  4.320 1.260 7.080 1.420 ;
        RECT  6.440 1.120 7.080 1.420 ;
        RECT  4.320 1.120 4.960 1.420 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.538  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.300 0.800 7.500 1.280 ;
        RECT  3.860 0.800 7.500 0.960 ;
        RECT  5.360 0.800 6.000 1.100 ;
        RECT  3.860 0.800 4.020 1.320 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.461  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 0.800 3.500 1.280 ;
        RECT  0.240 0.800 3.500 0.960 ;
        RECT  1.600 0.800 1.880 1.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.461  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.260 3.080 1.420 ;
        RECT  2.440 1.120 3.080 1.420 ;
        RECT  0.100 1.240 1.400 1.420 ;
        RECT  0.760 1.120 1.400 1.420 ;
        RECT  0.100 1.240 0.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.888  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.940 1.580 7.900 1.740 ;
        RECT  7.700 0.480 7.900 1.740 ;
        RECT  0.860 0.480 7.900 0.640 ;
        RECT  0.860 0.310 1.060 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  2.620 1.900 2.900 2.540 ;
        RECT  0.940 1.900 1.220 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.500 -0.140 7.780 0.320 ;
        RECT  5.380 -0.140 6.020 0.320 ;
        RECT  3.620 -0.140 3.900 0.320 ;
        RECT  2.500 -0.140 2.780 0.320 ;
        RECT  1.380 -0.140 1.660 0.320 ;
        RECT  0.340 -0.140 0.540 0.590 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.600 1.580 3.740 1.740 ;
        RECT  3.460 1.540 3.740 2.060 ;
        RECT  1.820 1.580 2.020 1.930 ;
        RECT  0.600 1.580 0.760 1.960 ;
        RECT  0.140 1.800 0.760 1.960 ;
        RECT  3.460 1.900 7.900 2.060 ;
        RECT  0.140 1.800 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END AOI211M8HM

MACRO AOI211M4HM
    CLASS CORE ;
    FOREIGN AOI211M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.269  LAYER ME1  ;
        ANTENNAGATEAREA 0.269  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.722  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.120 3.100 1.320 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.640 1.120 3.280 1.370 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.269  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.560 0.800 3.900 1.280 ;
        RECT  2.180 0.800 3.900 0.960 ;
        RECT  2.180 0.800 2.340 1.320 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.660 0.800 1.900 1.280 ;
        RECT  0.240 0.800 1.900 0.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 1.440 1.280 ;
        RECT  0.100 1.120 0.300 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.260 1.580 4.300 1.740 ;
        RECT  4.100 0.480 4.300 1.740 ;
        RECT  1.420 0.480 4.300 0.640 ;
        RECT  1.420 0.360 1.620 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  0.980 1.840 1.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.700 -0.140 3.980 0.320 ;
        RECT  1.940 -0.140 2.220 0.320 ;
        RECT  0.900 -0.140 1.100 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.600 1.520 2.060 1.680 ;
        RECT  1.780 1.520 2.060 2.060 ;
        RECT  0.600 1.520 0.760 1.960 ;
        RECT  0.140 1.800 0.760 1.960 ;
        RECT  1.780 1.900 4.140 2.060 ;
        RECT  0.140 1.800 0.340 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AOI211M4HM

MACRO AOI211M2HM
    CLASS CORE ;
    FOREIGN AOI211M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.300 1.510 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.840 1.540 1.420 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.000 1.100 1.670 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.480 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.542  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.640 0.480 2.300 0.680 ;
        RECT  1.460 1.580 1.900 1.740 ;
        RECT  1.700 0.480 1.900 1.740 ;
        RECT  0.640 0.480 0.840 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  0.180 1.480 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.980 1.900 2.300 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI211M2HM

MACRO AOI211M1HM
    CLASS CORE ;
    FOREIGN AOI211M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.300 1.510 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.098  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.840 1.540 1.420 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.970 1.100 1.640 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.470 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.423  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.620 0.480 2.300 0.680 ;
        RECT  1.460 1.580 1.900 1.740 ;
        RECT  1.700 0.480 1.900 1.740 ;
        RECT  0.620 0.480 0.900 0.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  0.300 1.800 0.500 2.540 ;
        RECT  0.140 1.800 0.500 2.000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.320 ;
        RECT  0.100 -0.140 0.380 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.980 1.800 1.260 2.100 ;
        RECT  2.080 1.740 2.280 2.100 ;
        RECT  0.980 1.900 2.280 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI211M1HM

MACRO AOI211M0HM
    CLASS CORE ;
    FOREIGN AOI211M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.300 1.510 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.079  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.840 1.540 1.420 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 1.000 1.100 1.670 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.065  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.480 1.280 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.358  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 0.480 2.300 0.680 ;
        RECT  1.460 1.580 1.900 1.780 ;
        RECT  1.700 0.480 1.900 1.780 ;
        RECT  0.660 0.480 0.860 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.400 2.540 ;
        RECT  0.180 1.490 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.400 0.140 ;
        RECT  1.140 -0.140 1.420 0.320 ;
        RECT  0.100 -0.140 0.380 0.320 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 2.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.400 1.140 ;
    END
END AOI211M0HM

MACRO AO33M8HM
    CLASS CORE ;
    FOREIGN AO33M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.695  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.120 4.700 1.320 ;
        LAYER ME2 ;
        RECT  4.500 1.040 4.700 1.560 ;
        LAYER ME1 ;
        RECT  4.180 1.020 4.760 1.410 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.555  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.120 5.900 1.320 ;
        LAYER ME2 ;
        RECT  5.700 1.040 5.900 1.560 ;
        LAYER ME1 ;
        RECT  5.360 1.120 6.000 1.370 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.027  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.120 3.100 1.320 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.400 1.040 3.240 1.360 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.320 0.800 6.700 1.280 ;
        RECT  4.920 0.800 6.700 0.960 ;
        RECT  4.920 0.800 5.080 1.320 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.880 0.800 2.040 1.360 ;
        RECT  0.460 0.800 2.040 0.960 ;
        RECT  0.460 0.800 0.700 1.360 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.700 1.540 9.100 2.100 ;
        RECT  8.900 0.370 9.100 2.100 ;
        RECT  7.700 0.660 9.100 0.860 ;
        RECT  8.760 0.370 9.100 0.860 ;
        RECT  7.660 1.540 9.100 1.740 ;
        RECT  7.660 1.540 7.940 2.100 ;
        RECT  7.700 0.390 7.900 0.860 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.555  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.120 1.500 1.320 ;
        LAYER ME2 ;
        RECT  1.300 1.040 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 1.120 1.600 1.370 ;
        END
    END B3
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  9.260 1.840 9.460 2.540 ;
        RECT  8.180 1.900 8.460 2.540 ;
        RECT  7.140 1.900 7.420 2.540 ;
        RECT  2.780 1.860 3.060 2.540 ;
        RECT  1.660 1.860 1.940 2.540 ;
        RECT  0.620 1.860 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  9.260 -0.140 9.460 0.560 ;
        RECT  8.180 -0.140 8.460 0.500 ;
        RECT  7.180 -0.140 7.380 0.670 ;
        RECT  5.580 -0.140 5.860 0.320 ;
        RECT  1.100 -0.140 1.380 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.020 0.300 3.380 0.460 ;
        RECT  3.100 0.300 3.380 0.520 ;
        RECT  2.020 0.300 2.220 0.640 ;
        RECT  0.180 0.480 2.220 0.640 ;
        RECT  3.580 0.300 5.000 0.460 ;
        RECT  4.620 0.300 5.000 0.640 ;
        RECT  3.580 0.300 3.860 0.520 ;
        RECT  4.620 0.480 6.780 0.640 ;
        RECT  0.100 1.540 3.580 1.700 ;
        RECT  3.340 1.540 3.580 2.100 ;
        RECT  0.100 1.540 0.380 2.100 ;
        RECT  1.140 1.540 1.420 2.100 ;
        RECT  2.180 1.540 2.460 2.100 ;
        RECT  3.340 1.900 6.900 2.100 ;
        RECT  2.540 0.620 2.820 0.860 ;
        RECT  4.140 0.620 4.420 0.860 ;
        RECT  2.540 0.700 4.420 0.860 ;
        RECT  7.340 1.040 8.700 1.240 ;
        RECT  3.740 0.700 3.900 1.740 ;
        RECT  7.340 1.040 7.500 1.740 ;
        RECT  3.740 1.580 7.500 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
    END
END AO33M8HM

MACRO AO33M4HM
    CLASS CORE ;
    FOREIGN AO33M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.866  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.100 3.500 1.300 ;
        LAYER ME2 ;
        RECT  3.300 1.020 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.000 1.040 3.500 1.360 ;
        END
    END B3
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 0.820 1.900 1.360 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.800 1.100 1.360 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.280 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.820 2.300 1.360 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.820 2.740 1.360 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 1.540 4.700 1.740 ;
        RECT  4.500 0.660 4.700 1.740 ;
        RECT  4.000 0.660 4.700 0.860 ;
        RECT  4.000 0.300 4.200 0.860 ;
        RECT  3.900 1.540 4.180 2.100 ;
        RECT  3.900 0.300 4.200 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.420 1.900 4.700 2.540 ;
        RECT  3.300 1.540 3.580 2.540 ;
        RECT  2.180 1.840 2.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.420 -0.140 4.700 0.500 ;
        RECT  3.280 -0.140 3.560 0.500 ;
        RECT  0.260 -0.140 0.460 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.660 1.520 2.980 1.680 ;
        RECT  0.620 1.840 0.900 2.100 ;
        RECT  1.660 1.520 1.940 2.100 ;
        RECT  0.620 1.940 1.940 2.100 ;
        RECT  2.700 1.520 2.980 2.100 ;
        RECT  1.260 0.360 3.120 0.520 ;
        RECT  2.960 0.360 3.120 0.820 ;
        RECT  2.960 0.660 3.820 0.820 ;
        RECT  3.660 0.660 3.820 1.300 ;
        RECT  3.660 1.020 4.320 1.300 ;
        RECT  0.100 1.520 1.420 1.680 ;
        RECT  1.260 0.360 1.420 1.780 ;
        RECT  1.140 1.520 1.420 1.780 ;
        RECT  0.100 1.520 0.380 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO33M4HM

MACRO AO33M2HM
    CLASS CORE ;
    FOREIGN AO33M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.800 2.340 1.360 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 0.840 1.900 1.360 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.100 1.070 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.280 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.800 2.820 1.360 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.580 1.560 ;
        RECT  3.080 1.040 3.580 1.360 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.390 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.440 1.730 3.640 2.540 ;
        RECT  2.260 1.840 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.380 -0.140 3.660 0.500 ;
        RECT  0.260 -0.140 0.460 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.800 1.520 3.020 1.680 ;
        RECT  0.620 1.840 0.900 2.100 ;
        RECT  2.820 1.520 3.020 2.010 ;
        RECT  1.800 1.520 1.960 2.100 ;
        RECT  0.620 1.940 1.960 2.100 ;
        RECT  1.260 0.360 3.220 0.520 ;
        RECT  3.060 0.360 3.220 0.820 ;
        RECT  3.060 0.660 3.900 0.820 ;
        RECT  3.740 0.660 3.900 1.320 ;
        RECT  0.140 1.520 1.460 1.680 ;
        RECT  1.260 0.360 1.460 1.780 ;
        RECT  1.100 1.520 1.460 1.780 ;
        RECT  0.140 1.520 0.340 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO33M2HM

MACRO AO33M1HM
    CLASS CORE ;
    FOREIGN AO33M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.750 2.340 1.320 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 0.840 1.900 1.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.100 1.120 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.280 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.800 2.820 1.320 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.580 1.560 ;
        RECT  3.080 1.040 3.580 1.360 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.390 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.440 1.730 3.640 2.540 ;
        RECT  2.260 1.840 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.380 -0.140 3.660 0.500 ;
        RECT  0.260 -0.140 0.460 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.800 1.520 3.020 1.680 ;
        RECT  0.620 1.840 0.900 2.100 ;
        RECT  2.820 1.520 3.020 2.010 ;
        RECT  1.800 1.520 1.960 2.100 ;
        RECT  0.620 1.940 1.960 2.100 ;
        RECT  1.260 0.360 3.220 0.520 ;
        RECT  3.060 0.360 3.220 0.820 ;
        RECT  3.060 0.660 3.900 0.820 ;
        RECT  3.740 0.660 3.900 1.320 ;
        RECT  0.140 1.520 1.460 1.680 ;
        RECT  1.260 0.360 1.460 1.780 ;
        RECT  1.180 1.520 1.460 1.780 ;
        RECT  0.140 1.520 0.340 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO33M1HM

MACRO AO33M0HM
    CLASS CORE ;
    FOREIGN AO33M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.750 2.340 1.360 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.620 0.840 1.900 1.360 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.100 1.160 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.360 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.800 2.820 1.360 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.082  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.300 1.040 3.580 1.560 ;
        RECT  3.080 1.040 3.580 1.360 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.310 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.440 1.730 3.640 2.540 ;
        RECT  2.260 1.840 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.380 -0.140 3.660 0.500 ;
        RECT  0.260 -0.140 0.460 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.800 1.520 3.020 1.680 ;
        RECT  0.620 1.840 0.900 2.100 ;
        RECT  2.820 1.520 3.020 2.010 ;
        RECT  1.800 1.520 1.960 2.100 ;
        RECT  0.620 1.940 1.960 2.100 ;
        RECT  1.260 0.360 3.220 0.520 ;
        RECT  3.060 0.360 3.220 0.820 ;
        RECT  3.060 0.660 3.900 0.820 ;
        RECT  3.740 0.660 3.900 1.320 ;
        RECT  0.140 1.520 1.460 1.680 ;
        RECT  1.260 0.360 1.460 1.780 ;
        RECT  1.180 1.520 1.460 1.780 ;
        RECT  0.140 1.520 0.340 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO33M0HM

MACRO AO32M8HM
    CLASS CORE ;
    FOREIGN AO32M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.712  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.160 2.700 1.360 ;
        LAYER ME2 ;
        RECT  2.500 1.080 2.700 1.600 ;
        LAYER ME1 ;
        RECT  2.380 1.080 3.060 1.380 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        ANTENNAGATEAREA 0.298  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.555  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.500 1.160 4.700 1.360 ;
        LAYER ME2 ;
        RECT  4.500 1.080 4.700 1.600 ;
        LAYER ME1 ;
        RECT  4.240 1.120 4.880 1.370 ;
        END
    END A3
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.600  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.160 1.500 1.360 ;
        LAYER ME2 ;
        RECT  1.300 1.080 1.500 1.600 ;
        LAYER ME1 ;
        RECT  1.000 1.120 1.640 1.370 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.298  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.220 0.800 5.380 1.360 ;
        RECT  3.700 0.800 5.380 0.960 ;
        RECT  3.700 0.800 3.940 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.800 2.060 1.360 ;
        RECT  0.460 0.800 2.060 0.960 ;
        RECT  0.460 0.800 0.700 1.360 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.500 1.540 7.900 2.080 ;
        RECT  7.700 0.350 7.900 2.080 ;
        RECT  6.500 0.660 7.900 0.860 ;
        RECT  7.560 0.350 7.900 0.860 ;
        RECT  6.460 1.540 7.900 1.740 ;
        RECT  6.460 1.540 6.740 2.080 ;
        RECT  6.500 0.390 6.700 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  8.060 1.800 8.260 2.540 ;
        RECT  6.980 1.900 7.260 2.540 ;
        RECT  5.980 1.450 6.180 2.540 ;
        RECT  1.700 1.860 1.980 2.540 ;
        RECT  0.660 1.860 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  8.060 -0.140 8.260 0.600 ;
        RECT  6.980 -0.140 7.260 0.500 ;
        RECT  5.980 -0.140 6.180 0.670 ;
        RECT  4.460 -0.140 4.740 0.320 ;
        RECT  1.140 -0.140 1.420 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.540 0.300 3.880 0.460 ;
        RECT  3.580 0.300 3.880 0.640 ;
        RECT  2.540 0.300 2.820 0.540 ;
        RECT  3.580 0.480 5.660 0.640 ;
        RECT  0.140 1.540 2.500 1.700 ;
        RECT  2.220 1.540 2.500 2.060 ;
        RECT  2.220 1.900 5.780 2.060 ;
        RECT  0.140 1.540 0.420 2.080 ;
        RECT  1.180 1.540 1.460 2.080 ;
        RECT  0.220 0.480 2.380 0.640 ;
        RECT  2.220 0.480 2.380 0.920 ;
        RECT  3.060 0.620 3.380 0.920 ;
        RECT  2.220 0.760 3.380 0.920 ;
        RECT  5.660 1.040 7.500 1.240 ;
        RECT  3.220 0.620 3.380 1.740 ;
        RECT  5.660 1.040 5.820 1.740 ;
        RECT  2.700 1.580 5.820 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
    END
END AO32M8HM

MACRO AO32M4HM
    CLASS CORE ;
    FOREIGN AO32M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.510  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.120 3.100 1.320 ;
        LAYER ME2 ;
        RECT  2.900 1.040 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.040 3.160 1.360 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 0.840 1.900 1.360 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.440 1.100 1.260 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.280 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.300 1.380 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 1.540 4.700 1.740 ;
        RECT  4.500 0.660 4.700 1.740 ;
        RECT  3.940 0.660 4.700 0.840 ;
        RECT  3.900 1.540 4.180 2.080 ;
        RECT  3.940 0.390 4.140 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.420 1.900 4.700 2.540 ;
        RECT  3.420 1.450 3.620 2.540 ;
        RECT  2.180 1.860 2.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.420 -0.140 4.700 0.500 ;
        RECT  3.380 -0.140 3.660 0.500 ;
        RECT  2.780 -0.140 3.060 0.500 ;
        RECT  0.260 -0.140 0.460 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.660 1.540 2.980 1.700 ;
        RECT  0.620 1.860 0.900 2.080 ;
        RECT  1.660 1.540 1.940 2.080 ;
        RECT  0.620 1.920 1.940 2.080 ;
        RECT  2.700 1.540 2.980 2.100 ;
        RECT  1.260 0.360 2.620 0.520 ;
        RECT  2.460 0.360 2.620 0.820 ;
        RECT  2.460 0.660 3.750 0.820 ;
        RECT  3.590 0.660 3.750 1.280 ;
        RECT  3.590 1.000 4.320 1.280 ;
        RECT  0.100 1.540 1.420 1.700 ;
        RECT  1.260 0.360 1.420 1.760 ;
        RECT  1.100 1.540 1.420 1.760 ;
        RECT  0.100 1.540 0.380 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO32M4HM

MACRO AO32M2HM
    CLASS CORE ;
    FOREIGN AO32M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.718  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.040 3.100 1.240 ;
        LAYER ME2 ;
        RECT  2.900 0.960 3.100 1.650 ;
        LAYER ME1 ;
        RECT  2.500 0.980 3.160 1.270 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 0.840 1.900 1.270 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.430 1.100 1.080 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.350 0.840 0.700 1.270 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.300 1.270 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.390 3.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.100 2.000 3.300 2.540 ;
        RECT  2.180 1.750 2.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.900 -0.140 3.180 0.500 ;
        RECT  0.260 -0.140 0.460 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.720 1.430 3.060 1.590 ;
        RECT  2.750 1.430 3.060 1.780 ;
        RECT  0.620 1.750 0.900 2.100 ;
        RECT  1.720 1.430 1.880 2.100 ;
        RECT  0.620 1.940 1.880 2.100 ;
        RECT  1.260 0.360 2.740 0.520 ;
        RECT  2.580 0.360 2.740 0.820 ;
        RECT  2.580 0.660 3.500 0.820 ;
        RECT  3.340 0.660 3.500 1.310 ;
        RECT  0.140 1.430 1.420 1.590 ;
        RECT  1.260 0.360 1.420 1.780 ;
        RECT  1.140 1.430 1.420 1.780 ;
        RECT  0.140 1.430 0.340 1.870 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END AO32M2HM

MACRO AO32M1HM
    CLASS CORE ;
    FOREIGN AO32M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.718  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.040 3.100 1.240 ;
        LAYER ME2 ;
        RECT  2.900 0.960 3.100 1.630 ;
        LAYER ME1 ;
        RECT  2.500 0.980 3.160 1.270 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 0.840 1.900 1.270 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.430 1.100 1.270 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 0.840 0.700 1.270 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.300 1.270 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.390 3.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.100 2.000 3.300 2.540 ;
        RECT  2.180 1.750 2.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.900 -0.140 3.180 0.500 ;
        RECT  0.260 -0.140 0.460 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.720 1.430 3.060 1.590 ;
        RECT  2.750 1.430 3.060 1.780 ;
        RECT  0.620 1.750 0.900 2.100 ;
        RECT  1.720 1.430 1.880 2.100 ;
        RECT  0.620 1.940 1.880 2.100 ;
        RECT  1.260 0.360 2.740 0.520 ;
        RECT  2.580 0.360 2.740 0.820 ;
        RECT  2.580 0.660 3.500 0.820 ;
        RECT  3.340 0.660 3.500 1.310 ;
        RECT  0.140 1.430 1.420 1.590 ;
        RECT  1.260 0.360 1.420 1.780 ;
        RECT  1.140 1.430 1.420 1.780 ;
        RECT  0.140 1.430 0.340 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END AO32M1HM

MACRO AO32M0HM
    CLASS CORE ;
    FOREIGN AO32M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.718  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.900 1.040 3.100 1.240 ;
        LAYER ME2 ;
        RECT  2.900 0.960 3.100 1.560 ;
        LAYER ME1 ;
        RECT  2.500 0.980 3.160 1.270 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.580 0.840 1.900 1.270 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.430 1.100 1.130 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.091  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.270 ;
        END
    END A3
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.100 0.750 2.300 1.270 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.680 0.310 3.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.100 2.000 3.300 2.540 ;
        RECT  2.180 1.750 2.460 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  2.900 -0.140 3.180 0.500 ;
        RECT  0.260 -0.140 0.460 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.720 1.430 3.060 1.590 ;
        RECT  2.750 1.430 3.060 1.780 ;
        RECT  0.620 1.750 0.900 2.100 ;
        RECT  1.720 1.430 1.880 2.100 ;
        RECT  0.620 1.940 1.880 2.100 ;
        RECT  1.260 0.360 2.740 0.520 ;
        RECT  2.580 0.360 2.740 0.820 ;
        RECT  2.580 0.660 3.500 0.820 ;
        RECT  3.340 0.660 3.500 1.310 ;
        RECT  0.140 1.430 1.420 1.590 ;
        RECT  1.260 0.360 1.420 1.780 ;
        RECT  1.140 1.430 1.420 1.780 ;
        RECT  0.140 1.430 0.340 1.970 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END AO32M0HM

MACRO AO31M8HM
    CLASS CORE ;
    FOREIGN AO31M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.295  LAYER ME2  ;
        ANTENNAGATEAREA 0.295  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.691  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.120 3.500 1.320 ;
        LAYER ME2 ;
        RECT  3.300 1.040 3.500 1.560 ;
        LAYER ME1 ;
        RECT  2.920 1.040 3.560 1.360 ;
        END
    END A1
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.295  LAYER ME1  ;
        ANTENNAGATEAREA 0.295  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.568  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.170 1.500 1.370 ;
        LAYER ME2 ;
        RECT  1.300 1.030 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.000 1.120 1.640 1.370 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.295  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.920 0.800 2.080 1.320 ;
        RECT  0.500 0.800 2.080 0.960 ;
        RECT  0.500 0.800 0.700 1.360 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.700 1.540 7.100 2.080 ;
        RECT  6.900 0.390 7.100 2.080 ;
        RECT  5.700 0.660 7.100 0.860 ;
        RECT  6.700 0.390 7.100 0.860 ;
        RECT  5.660 1.540 7.100 1.740 ;
        RECT  5.660 1.540 5.940 2.080 ;
        RECT  5.700 0.390 5.900 0.860 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.250  LAYER ME1  ;
        ANTENNAGATEAREA 0.250  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.000  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.120 4.300 1.320 ;
        LAYER ME2 ;
        RECT  4.100 1.040 4.300 1.560 ;
        LAYER ME1 ;
        RECT  3.960 1.040 4.600 1.360 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.600 2.540 ;
        RECT  7.260 1.480 7.460 2.540 ;
        RECT  6.180 1.900 6.460 2.540 ;
        RECT  5.180 1.450 5.380 2.540 ;
        RECT  4.140 1.860 4.420 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.600 0.140 ;
        RECT  7.260 -0.140 7.460 0.600 ;
        RECT  6.180 -0.140 6.460 0.500 ;
        RECT  5.140 -0.140 5.420 0.500 ;
        RECT  4.140 -0.140 4.420 0.500 ;
        RECT  1.140 -0.140 1.440 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.070 0.300 3.380 0.460 ;
        RECT  3.100 0.300 3.380 0.500 ;
        RECT  2.070 0.300 2.340 0.640 ;
        RECT  0.220 0.480 2.340 0.640 ;
        RECT  3.620 1.540 4.940 1.700 ;
        RECT  0.140 1.540 0.420 2.060 ;
        RECT  3.620 1.540 3.900 2.060 ;
        RECT  0.140 1.900 3.900 2.060 ;
        RECT  4.660 1.540 4.940 2.080 ;
        RECT  2.540 0.620 2.860 0.820 ;
        RECT  3.660 0.330 3.860 0.820 ;
        RECT  4.700 0.310 4.900 0.820 ;
        RECT  2.540 0.660 5.480 0.820 ;
        RECT  5.320 0.660 5.480 1.240 ;
        RECT  5.320 1.040 6.620 1.240 ;
        RECT  2.540 0.620 2.760 1.740 ;
        RECT  0.620 1.580 3.420 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.600 1.140 ;
    END
END AO31M8HM

MACRO AO31M4HM
    CLASS CORE ;
    FOREIGN AO31M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        ANTENNAGATEAREA 0.127  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.434  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.120 2.300 1.320 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.800 1.040 2.300 1.380 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.260 0.840 1.540 1.420 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.440 1.100 1.280 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.200 0.840 0.700 1.360 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.800 1.540 3.500 1.740 ;
        RECT  3.300 0.660 3.500 1.740 ;
        RECT  2.800 0.660 3.500 0.860 ;
        RECT  2.700 1.900 3.000 2.100 ;
        RECT  2.800 1.540 3.000 2.100 ;
        RECT  2.800 0.300 3.000 0.860 ;
        RECT  2.700 0.300 3.000 0.500 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.180 -0.140 2.460 0.500 ;
        RECT  0.220 -0.140 0.420 0.640 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.620 1.900 1.940 2.100 ;
        RECT  1.700 0.300 1.860 0.820 ;
        RECT  1.700 0.660 2.620 0.820 ;
        RECT  2.460 1.040 3.120 1.320 ;
        RECT  2.460 0.660 2.620 1.740 ;
        RECT  0.140 1.580 2.620 1.740 ;
        RECT  0.140 1.580 0.340 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AO31M4HM

MACRO AO31M2HM
    CLASS CORE ;
    FOREIGN AO31M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.120 2.300 1.320 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.960 2.380 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.640 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.760 1.140 1.280 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.280 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.390 3.100 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.240 -0.140 2.520 0.480 ;
        RECT  0.300 -0.140 0.500 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.900 0.940 2.100 ;
        RECT  1.700 1.900 1.980 2.100 ;
        RECT  0.660 1.940 1.980 2.100 ;
        RECT  1.620 0.380 2.000 0.580 ;
        RECT  1.840 0.380 2.000 0.800 ;
        RECT  1.840 0.640 2.700 0.800 ;
        RECT  2.540 0.640 2.700 1.740 ;
        RECT  0.180 1.580 2.700 1.740 ;
        RECT  1.140 1.580 1.500 1.780 ;
        RECT  0.180 1.580 0.380 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO31M2HM

MACRO AO31M1HM
    CLASS CORE ;
    FOREIGN AO31M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.120 2.300 1.320 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.960 2.380 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.640 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.770 1.140 1.280 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.480 0.770 0.700 1.280 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.390 3.100 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.240 -0.140 2.520 0.480 ;
        RECT  0.300 -0.140 0.500 0.610 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.900 0.940 2.100 ;
        RECT  1.700 1.900 1.980 2.100 ;
        RECT  0.660 1.940 1.980 2.100 ;
        RECT  1.620 0.380 2.040 0.580 ;
        RECT  1.880 0.380 2.040 0.800 ;
        RECT  1.880 0.640 2.700 0.800 ;
        RECT  2.540 0.640 2.700 1.740 ;
        RECT  0.180 1.580 2.700 1.740 ;
        RECT  1.140 1.580 1.500 1.780 ;
        RECT  0.180 1.580 0.380 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO31M1HM

MACRO AO31M0HM
    CLASS CORE ;
    FOREIGN AO31M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.120 2.300 1.320 ;
        LAYER ME2 ;
        RECT  2.100 1.040 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.960 2.380 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.640 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.140 1.280 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.280 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.880 0.310 3.100 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.260 1.900 2.540 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.240 -0.140 2.520 0.480 ;
        RECT  0.300 -0.140 0.500 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 1.900 0.940 2.100 ;
        RECT  1.700 1.900 1.980 2.100 ;
        RECT  0.660 1.940 1.980 2.100 ;
        RECT  1.620 0.380 2.030 0.580 ;
        RECT  1.870 0.380 2.030 0.800 ;
        RECT  1.870 0.640 2.700 0.800 ;
        RECT  2.540 0.640 2.700 1.740 ;
        RECT  0.180 1.580 2.700 1.740 ;
        RECT  1.140 1.580 1.500 1.780 ;
        RECT  0.180 1.580 0.380 1.960 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO31M0HM

MACRO AO22M8HM
    CLASS CORE ;
    FOREIGN AO22M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.960 0.850 3.640 1.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.620 1.260 4.140 1.420 ;
        RECT  3.980 0.850 4.140 1.420 ;
        RECT  2.620 0.850 2.780 1.420 ;
        RECT  2.440 0.850 2.780 1.230 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.110 0.850 1.720 1.100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.260 2.060 1.420 ;
        RECT  1.900 0.930 2.060 1.420 ;
        RECT  0.500 0.840 0.700 1.420 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 0.370 6.540 2.100 ;
        RECT  5.260 1.520 6.540 1.720 ;
        RECT  6.100 0.660 6.540 1.720 ;
        RECT  5.300 0.660 6.540 0.840 ;
        RECT  5.260 1.520 5.500 2.100 ;
        RECT  5.300 0.370 5.500 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.860 1.460 7.060 2.540 ;
        RECT  5.780 1.880 6.060 2.540 ;
        RECT  4.740 1.430 5.020 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.860 -0.140 7.060 0.720 ;
        RECT  5.780 -0.140 6.060 0.500 ;
        RECT  4.740 -0.140 4.940 0.690 ;
        RECT  4.140 -0.140 4.420 0.340 ;
        RECT  2.300 -0.140 2.580 0.340 ;
        RECT  0.220 -0.140 0.500 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.130 1.580 2.420 1.740 ;
        RECT  2.220 1.580 2.420 2.060 ;
        RECT  1.180 1.580 1.380 1.960 ;
        RECT  0.130 1.580 0.340 1.970 ;
        RECT  2.220 1.900 4.580 2.060 ;
        RECT  1.080 0.530 4.500 0.690 ;
        RECT  4.300 1.040 5.790 1.240 ;
        RECT  4.300 0.530 4.500 1.740 ;
        RECT  2.660 1.580 4.500 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END AO22M8HM

MACRO AO22M4HM
    CLASS CORE ;
    FOREIGN AO22M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.460 0.980 2.700 1.650 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.020 1.000 1.500 1.280 ;
        RECT  1.300 0.840 1.500 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.280 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.040 2.180 1.240 ;
        RECT  1.700 1.040 1.900 1.560 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.140 1.460 3.900 1.660 ;
        RECT  3.700 0.700 3.900 1.660 ;
        RECT  3.260 0.700 3.900 0.900 ;
        RECT  3.260 0.300 3.460 0.900 ;
        RECT  3.140 1.460 3.340 2.100 ;
        RECT  3.100 0.300 3.460 0.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.000 2.540 ;
        RECT  3.620 1.820 3.900 2.540 ;
        RECT  2.620 1.810 2.820 2.540 ;
        RECT  1.500 2.080 1.780 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.000 0.140 ;
        RECT  3.620 -0.140 3.900 0.540 ;
        RECT  2.580 -0.140 2.860 0.500 ;
        RECT  0.320 -0.140 0.520 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 1.440 1.360 1.920 ;
        RECT  1.000 1.760 2.280 1.920 ;
        RECT  0.100 1.880 1.160 2.040 ;
        RECT  2.120 1.460 2.280 2.100 ;
        RECT  0.680 0.440 2.360 0.600 ;
        RECT  2.200 0.440 2.360 0.820 ;
        RECT  2.200 0.660 3.060 0.820 ;
        RECT  2.900 0.660 3.060 1.220 ;
        RECT  2.900 1.060 3.380 1.220 ;
        RECT  0.680 0.440 0.840 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.000 1.140 ;
    END
END AO22M4HM

MACRO AO22M2HM
    CLASS CORE ;
    FOREIGN AO22M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.755  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.140 1.140 2.340 1.340 ;
        LAYER ME2 ;
        RECT  2.100 0.850 2.340 1.570 ;
        LAYER ME1 ;
        RECT  2.140 1.000 2.490 1.440 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.360 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.320 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.370 3.500 2.100 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.700 -0.140 2.980 0.520 ;
        RECT  2.020 -0.140 2.300 0.500 ;
        RECT  0.220 -0.140 0.420 0.580 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.700 1.530 2.980 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.160 1.580 1.360 1.740 ;
        RECT  1.200 1.580 1.360 2.060 ;
        RECT  2.220 1.690 2.500 2.060 ;
        RECT  1.200 1.900 2.500 2.060 ;
        RECT  0.160 1.580 0.320 2.100 ;
        RECT  1.040 0.340 1.860 0.500 ;
        RECT  1.700 0.680 3.100 0.840 ;
        RECT  2.940 0.680 3.100 1.370 ;
        RECT  1.700 0.340 1.860 1.740 ;
        RECT  1.700 1.520 1.980 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AO22M2HM

MACRO AO22M1HM
    CLASS CORE ;
    FOREIGN AO22M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.755  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.140 1.140 2.340 1.340 ;
        LAYER ME2 ;
        RECT  2.100 0.850 2.340 1.570 ;
        LAYER ME1 ;
        RECT  2.140 1.000 2.490 1.440 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.360 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.840 0.700 1.320 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.370 3.500 1.960 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.700 -0.140 2.980 0.520 ;
        RECT  2.020 -0.140 2.300 0.500 ;
        RECT  0.220 -0.140 0.420 0.580 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.740 1.530 2.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.160 1.580 1.360 1.740 ;
        RECT  1.200 1.580 1.360 2.060 ;
        RECT  2.220 1.690 2.500 2.060 ;
        RECT  1.200 1.900 2.500 2.060 ;
        RECT  0.160 1.580 0.320 2.100 ;
        RECT  1.040 0.340 1.860 0.500 ;
        RECT  1.700 0.680 3.100 0.840 ;
        RECT  2.940 0.680 3.100 1.370 ;
        RECT  1.700 0.340 1.860 1.740 ;
        RECT  1.700 1.520 1.980 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AO22M1HM

MACRO AO22M0HM
    CLASS CORE ;
    FOREIGN AO22M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.280 0.300 3.500 1.960 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.755  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.140 1.140 2.340 1.340 ;
        LAYER ME2 ;
        RECT  2.100 0.850 2.340 1.570 ;
        LAYER ME1 ;
        RECT  2.140 1.000 2.490 1.440 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.360 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.360 0.840 0.700 1.320 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.700 -0.140 2.980 0.520 ;
        RECT  2.020 -0.140 2.300 0.500 ;
        RECT  0.220 -0.140 0.420 0.580 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.740 1.530 2.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.160 1.580 1.360 1.740 ;
        RECT  1.200 1.580 1.360 2.060 ;
        RECT  2.220 1.690 2.500 2.060 ;
        RECT  1.200 1.900 2.500 2.060 ;
        RECT  0.160 1.580 0.320 2.100 ;
        RECT  1.040 0.340 1.860 0.500 ;
        RECT  1.700 0.680 3.100 0.840 ;
        RECT  2.940 0.680 3.100 1.370 ;
        RECT  1.700 0.340 1.860 1.740 ;
        RECT  1.700 1.520 1.980 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AO22M0HM

MACRO AO22B11M8HM
    CLASS CORE ;
    FOREIGN AO22B11M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.940 0.800 5.240 1.100 ;
        RECT  3.480 0.800 5.240 0.960 ;
        RECT  3.480 0.800 3.960 1.210 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.840 0.800 3.000 1.320 ;
        RECT  1.070 0.800 3.000 0.960 ;
        RECT  1.070 0.800 1.560 1.100 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.940 0.840 6.300 1.320 ;
        END
    END NA2
    PIN NB2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.400 ;
        END
    END NB2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.040 0.900 8.360 1.160 ;
        RECT  7.820 1.540 8.240 2.100 ;
        RECT  8.040 0.370 8.240 2.100 ;
        RECT  6.840 0.660 8.240 0.860 ;
        RECT  7.880 0.370 8.240 0.860 ;
        RECT  6.770 1.540 8.240 1.740 ;
        RECT  6.770 1.540 7.100 2.100 ;
        RECT  6.840 0.370 7.040 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.400 1.450 8.600 2.540 ;
        RECT  7.320 1.900 7.600 2.540 ;
        RECT  6.320 1.760 6.520 2.540 ;
        RECT  2.600 2.020 2.880 2.540 ;
        RECT  1.520 1.900 1.800 2.540 ;
        RECT  0.140 1.560 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.400 -0.140 8.600 0.650 ;
        RECT  7.320 -0.140 7.600 0.500 ;
        RECT  6.240 -0.140 6.520 0.320 ;
        RECT  4.120 -0.140 4.400 0.320 ;
        RECT  2.000 -0.140 2.280 0.320 ;
        RECT  0.140 -0.140 0.340 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.680 0.310 0.840 1.420 ;
        RECT  1.830 1.120 2.500 1.420 ;
        RECT  0.680 1.260 2.500 1.420 ;
        RECT  0.720 1.260 0.880 1.700 ;
        RECT  1.140 1.580 3.000 1.740 ;
        RECT  2.840 1.690 3.400 1.850 ;
        RECT  3.200 1.690 3.400 2.100 ;
        RECT  4.150 1.900 4.500 2.100 ;
        RECT  2.020 1.580 2.340 1.980 ;
        RECT  1.140 1.580 1.300 2.100 ;
        RECT  0.860 1.940 1.300 2.100 ;
        RECT  5.280 1.800 5.480 2.100 ;
        RECT  3.200 1.940 5.480 2.100 ;
        RECT  4.150 1.120 4.530 1.420 ;
        RECT  5.480 0.620 5.760 1.420 ;
        RECT  4.150 1.260 5.760 1.420 ;
        RECT  5.580 0.620 5.760 1.640 ;
        RECT  5.760 1.480 5.960 2.020 ;
        RECT  5.000 0.300 6.080 0.460 ;
        RECT  5.920 0.300 6.080 0.640 ;
        RECT  5.000 0.300 5.280 0.640 ;
        RECT  1.020 0.480 5.280 0.640 ;
        RECT  5.920 0.480 6.620 0.640 ;
        RECT  6.460 0.480 6.620 1.240 ;
        RECT  6.460 1.040 7.840 1.240 ;
        RECT  3.160 0.480 3.320 1.530 ;
        RECT  3.160 1.370 3.850 1.530 ;
        RECT  3.680 1.370 3.850 1.780 ;
        RECT  3.680 1.580 5.080 1.740 ;
        RECT  3.680 1.580 4.000 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.080 1.760 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.080 ;
        RECT  1.760 0.000 8.800 1.140 ;
    END
END AO22B11M8HM

MACRO AO22B11M4HM
    CLASS CORE ;
    FOREIGN AO22B11M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.507  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.080 1.900 1.280 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.700 0.980 2.040 1.340 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.722  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.400 1.140 2.600 1.340 ;
        LAYER ME2 ;
        RECT  2.400 0.840 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.200 1.080 2.700 1.340 ;
        END
    END A1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.960 1.120 4.360 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.690 1.540 5.500 1.740 ;
        RECT  5.300 0.680 5.500 1.740 ;
        RECT  4.840 0.680 5.500 0.880 ;
        RECT  4.840 0.410 5.040 0.880 ;
        RECT  4.660 0.410 5.040 0.640 ;
        END
    END Z
    PIN NB2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        ANTENNAGATEAREA 0.083  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.961  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.620 0.620 0.820 0.820 ;
        LAYER ME2 ;
        RECT  0.500 0.440 0.820 1.160 ;
        LAYER ME1 ;
        RECT  0.520 0.480 0.860 0.930 ;
        END
    END NB2
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.600 2.540 ;
        RECT  5.220 1.900 5.500 2.540 ;
        RECT  4.180 1.900 4.460 2.540 ;
        RECT  1.540 1.900 1.820 2.540 ;
        RECT  0.660 2.080 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.600 0.140 ;
        RECT  5.220 -0.140 5.500 0.520 ;
        RECT  4.240 -0.140 4.440 0.640 ;
        RECT  1.980 -0.140 2.260 0.460 ;
        RECT  0.660 -0.140 0.940 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.100 1.520 1.300 ;
        RECT  0.100 0.310 0.320 2.100 ;
        RECT  0.980 1.500 2.350 1.700 ;
        RECT  2.080 1.500 2.350 2.100 ;
        RECT  2.080 1.880 3.390 2.100 ;
        RECT  3.480 0.620 3.760 1.340 ;
        RECT  3.600 0.620 3.760 2.030 ;
        RECT  3.600 1.830 3.940 2.030 ;
        RECT  2.860 0.300 4.080 0.460 ;
        RECT  1.020 0.620 3.090 0.780 ;
        RECT  3.920 0.300 4.080 0.960 ;
        RECT  3.920 0.800 4.680 0.960 ;
        RECT  4.520 0.800 4.680 1.320 ;
        RECT  4.520 1.040 5.120 1.320 ;
        RECT  2.860 0.300 3.090 1.720 ;
        RECT  2.550 1.560 3.090 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.600 1.140 ;
    END
END AO22B11M4HM

MACRO AO22B11M2HM
    CLASS CORE ;
    FOREIGN AO22B11M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.657  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.160 2.700 1.360 ;
        LAYER ME2 ;
        RECT  2.500 0.770 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.020 2.700 1.460 ;
        RECT  2.200 1.020 2.700 1.260 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 2.000 1.260 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.960 1.120 4.390 1.560 ;
        END
    END NA2
    PIN NB2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.300 ;
        END
    END NB2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.680 5.100 2.020 ;
        RECT  4.900 0.340 5.100 2.020 ;
        RECT  4.780 0.340 5.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  1.520 1.740 1.800 2.540 ;
        RECT  0.100 1.560 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.360 -0.140 4.560 0.640 ;
        RECT  2.820 -0.140 3.100 0.530 ;
        RECT  1.100 -0.140 1.300 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.540 0.340 0.880 0.540 ;
        RECT  0.720 0.980 1.520 1.180 ;
        RECT  0.720 0.340 0.880 1.700 ;
        RECT  1.120 1.420 2.320 1.580 ;
        RECT  2.100 1.420 2.320 2.100 ;
        RECT  1.120 1.420 1.280 2.100 ;
        RECT  0.900 1.940 1.280 2.100 ;
        RECT  3.200 1.590 3.420 2.100 ;
        RECT  2.100 1.940 3.420 2.100 ;
        RECT  3.600 0.620 3.880 0.910 ;
        RECT  3.180 1.010 3.760 1.290 ;
        RECT  3.600 0.620 3.760 2.030 ;
        RECT  3.600 1.830 3.940 2.030 ;
        RECT  3.280 0.300 4.200 0.460 ;
        RECT  1.870 0.370 2.550 0.530 ;
        RECT  2.390 0.370 2.550 0.860 ;
        RECT  4.040 0.300 4.200 0.960 ;
        RECT  3.280 0.300 3.440 0.850 ;
        RECT  2.390 0.690 3.440 0.850 ;
        RECT  2.390 0.690 3.020 0.860 ;
        RECT  4.040 0.800 4.740 0.960 ;
        RECT  4.580 0.800 4.740 1.390 ;
        RECT  2.860 0.690 3.020 1.780 ;
        RECT  2.520 1.620 3.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.010 1.210 2.400 ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.010 ;
        RECT  1.210 0.000 5.200 1.140 ;
    END
END AO22B11M2HM

MACRO AO22B11M1HM
    CLASS CORE ;
    FOREIGN AO22B11M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.657  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.160 2.700 1.360 ;
        LAYER ME2 ;
        RECT  2.500 0.770 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.020 2.700 1.460 ;
        RECT  2.200 1.020 2.700 1.260 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.840 2.000 1.260 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.960 1.120 4.390 1.560 ;
        END
    END NA2
    PIN NB2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.250 ;
        END
    END NB2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.680 5.100 2.020 ;
        RECT  4.900 0.340 5.100 2.020 ;
        RECT  4.780 0.340 5.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  1.520 1.740 1.800 2.540 ;
        RECT  0.100 1.560 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.360 -0.140 4.560 0.640 ;
        RECT  2.820 -0.140 3.100 0.530 ;
        RECT  1.100 -0.140 1.300 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.540 0.340 0.880 0.540 ;
        RECT  0.720 0.980 1.520 1.180 ;
        RECT  0.720 0.340 0.880 1.700 ;
        RECT  1.120 1.420 2.320 1.580 ;
        RECT  2.100 1.420 2.320 2.100 ;
        RECT  1.120 1.420 1.280 2.100 ;
        RECT  0.900 1.940 1.280 2.100 ;
        RECT  3.200 1.590 3.420 2.100 ;
        RECT  2.100 1.940 3.420 2.100 ;
        RECT  3.600 0.620 3.880 0.910 ;
        RECT  3.180 1.010 3.760 1.290 ;
        RECT  3.600 0.620 3.760 2.030 ;
        RECT  3.600 1.830 3.940 2.030 ;
        RECT  3.280 0.300 4.200 0.460 ;
        RECT  1.870 0.370 2.550 0.530 ;
        RECT  2.390 0.370 2.550 0.860 ;
        RECT  4.040 0.300 4.200 0.960 ;
        RECT  3.280 0.300 3.440 0.850 ;
        RECT  2.390 0.690 3.440 0.850 ;
        RECT  2.390 0.690 3.020 0.860 ;
        RECT  4.040 0.800 4.740 0.960 ;
        RECT  4.580 0.800 4.740 1.390 ;
        RECT  2.860 0.690 3.020 1.780 ;
        RECT  2.520 1.620 3.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.010 1.210 2.400 ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.010 ;
        RECT  1.210 0.000 5.200 1.140 ;
    END
END AO22B11M1HM

MACRO AO22B11M0HM
    CLASS CORE ;
    FOREIGN AO22B11M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.657  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.160 2.700 1.360 ;
        LAYER ME2 ;
        RECT  2.500 0.770 2.700 1.560 ;
        LAYER ME1 ;
        RECT  2.500 1.020 2.700 1.460 ;
        RECT  2.200 1.020 2.700 1.260 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.730 2.000 1.260 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.960 1.120 4.390 1.560 ;
        END
    END NA2
    PIN NB2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.500 1.300 ;
        END
    END NB2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.820 1.680 5.100 2.020 ;
        RECT  4.900 0.340 5.100 2.020 ;
        RECT  4.780 0.340 5.100 0.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.300 1.900 4.580 2.540 ;
        RECT  1.520 1.740 1.800 2.540 ;
        RECT  0.100 1.560 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.360 -0.140 4.560 0.640 ;
        RECT  2.820 -0.140 3.100 0.530 ;
        RECT  1.100 -0.140 1.300 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.540 0.340 0.880 0.540 ;
        RECT  0.720 0.940 1.520 1.220 ;
        RECT  0.720 0.340 0.880 1.700 ;
        RECT  1.120 1.420 2.320 1.580 ;
        RECT  2.100 1.420 2.320 2.100 ;
        RECT  1.120 1.420 1.280 2.100 ;
        RECT  0.900 1.940 1.280 2.100 ;
        RECT  3.200 1.590 3.420 2.100 ;
        RECT  2.100 1.940 3.420 2.100 ;
        RECT  3.600 0.620 3.880 0.910 ;
        RECT  3.180 1.010 3.760 1.290 ;
        RECT  3.600 0.620 3.760 2.030 ;
        RECT  3.600 1.830 3.940 2.030 ;
        RECT  3.280 0.300 4.200 0.460 ;
        RECT  1.870 0.370 2.550 0.530 ;
        RECT  2.390 0.370 2.550 0.860 ;
        RECT  4.040 0.300 4.200 0.960 ;
        RECT  3.280 0.300 3.440 0.850 ;
        RECT  2.390 0.690 3.440 0.850 ;
        RECT  2.390 0.690 3.020 0.860 ;
        RECT  4.040 0.800 4.740 0.960 ;
        RECT  4.580 0.800 4.740 1.390 ;
        RECT  2.860 0.690 3.020 1.780 ;
        RECT  2.520 1.620 3.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.010 1.210 2.400 ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.010 ;
        RECT  1.210 0.000 5.200 1.140 ;
    END
END AO22B11M0HM

MACRO AO22B10M8HM
    CLASS CORE ;
    FOREIGN AO22B10M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        ANTENNAGATEAREA 0.289  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.636  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.140 1.500 1.340 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.930 1.120 1.600 1.360 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.040 0.800 4.320 1.100 ;
        RECT  2.700 0.800 4.320 0.960 ;
        RECT  2.700 0.800 3.160 1.230 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.289  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.960 0.800 2.120 1.320 ;
        RECT  0.500 0.800 2.120 0.960 ;
        RECT  0.500 0.800 0.700 1.360 ;
        END
    END B1
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.101  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.180 0.840 5.500 1.320 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.080 1.540 7.500 2.100 ;
        RECT  7.300 0.370 7.500 2.100 ;
        RECT  6.100 0.660 7.500 0.860 ;
        RECT  7.140 0.370 7.500 0.860 ;
        RECT  6.030 1.540 7.500 1.740 ;
        RECT  6.030 1.540 6.360 2.100 ;
        RECT  6.100 0.370 6.300 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.660 1.450 7.860 2.540 ;
        RECT  6.580 1.900 6.860 2.540 ;
        RECT  5.580 1.720 5.780 2.540 ;
        RECT  1.700 2.000 1.920 2.540 ;
        RECT  0.620 1.880 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.660 -0.140 7.860 0.650 ;
        RECT  6.580 -0.140 6.860 0.500 ;
        RECT  5.500 -0.140 5.780 0.320 ;
        RECT  3.340 -0.140 3.620 0.320 ;
        RECT  1.180 -0.140 1.460 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.520 1.440 1.680 ;
        RECT  1.120 1.650 2.250 1.810 ;
        RECT  2.080 1.650 2.250 2.100 ;
        RECT  2.080 1.840 2.590 2.100 ;
        RECT  3.250 1.900 3.600 2.100 ;
        RECT  0.100 1.520 0.400 2.100 ;
        RECT  1.120 1.520 1.440 2.100 ;
        RECT  4.380 1.800 4.580 2.100 ;
        RECT  2.080 1.940 4.580 2.100 ;
        RECT  4.520 0.620 5.020 0.840 ;
        RECT  3.460 1.120 3.740 1.420 ;
        RECT  3.460 1.260 4.680 1.420 ;
        RECT  4.520 0.620 4.680 1.640 ;
        RECT  4.520 1.480 5.220 1.640 ;
        RECT  5.020 1.480 5.220 2.020 ;
        RECT  4.070 0.300 5.340 0.460 ;
        RECT  5.180 0.300 5.340 0.640 ;
        RECT  4.070 0.300 4.230 0.640 ;
        RECT  0.200 0.480 4.230 0.640 ;
        RECT  5.180 0.480 5.880 0.640 ;
        RECT  5.720 0.480 5.880 1.240 ;
        RECT  5.720 1.040 7.100 1.240 ;
        RECT  2.380 0.480 2.540 1.550 ;
        RECT  2.380 1.390 3.020 1.550 ;
        RECT  2.780 1.580 4.180 1.740 ;
        RECT  2.780 1.390 3.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
    END
END AO22B10M8HM

MACRO AO22B10M4HM
    CLASS CORE ;
    FOREIGN AO22B10M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        ANTENNAGATEAREA 0.145  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.937  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.080 2.300 1.280 ;
        LAYER ME2 ;
        RECT  2.100 0.990 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.940 2.460 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.340 1.280 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.980 1.320 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.180 1.140 3.560 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.870 1.540 4.700 1.740 ;
        RECT  4.500 0.680 4.700 1.740 ;
        RECT  4.080 0.680 4.700 0.880 ;
        RECT  4.080 0.300 4.240 0.880 ;
        RECT  3.870 1.540 4.190 2.100 ;
        RECT  3.850 0.300 4.240 0.510 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.420 1.900 4.700 2.540 ;
        RECT  3.420 1.810 3.620 2.540 ;
        RECT  0.660 1.950 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.420 -0.140 4.700 0.520 ;
        RECT  3.440 -0.140 3.640 0.560 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.630 1.440 1.790 ;
        RECT  1.280 1.630 1.440 2.100 ;
        RECT  0.100 1.440 0.390 2.100 ;
        RECT  2.260 1.520 2.540 2.100 ;
        RECT  1.280 1.940 2.540 2.100 ;
        RECT  1.740 0.620 2.960 0.780 ;
        RECT  1.740 0.620 1.900 1.000 ;
        RECT  1.460 0.840 1.740 1.150 ;
        RECT  2.800 0.620 2.960 1.990 ;
        RECT  2.800 1.770 3.100 1.990 ;
        RECT  1.420 0.300 3.280 0.460 ;
        RECT  0.100 0.420 0.400 0.680 ;
        RECT  1.420 0.300 1.580 0.680 ;
        RECT  0.100 0.480 1.580 0.680 ;
        RECT  3.120 0.300 3.280 0.880 ;
        RECT  3.120 0.720 3.880 0.880 ;
        RECT  3.720 0.720 3.880 1.320 ;
        RECT  1.140 0.480 1.300 1.470 ;
        RECT  3.720 1.040 4.320 1.320 ;
        RECT  1.140 1.310 1.860 1.470 ;
        RECT  1.700 1.310 1.860 1.780 ;
        RECT  1.700 1.620 2.060 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO22B10M4HM

MACRO AO22B10M2HM
    CLASS CORE ;
    FOREIGN AO22B10M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.935  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.080 2.300 1.280 ;
        LAYER ME2 ;
        RECT  2.100 0.990 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.940 2.460 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.340 1.280 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.980 1.320 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.180 1.140 3.560 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.870 1.540 4.300 2.100 ;
        RECT  4.100 0.300 4.300 2.100 ;
        RECT  3.850 0.300 4.300 0.510 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.420 1.810 3.620 2.540 ;
        RECT  0.660 1.950 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.440 -0.140 3.640 0.560 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.630 1.440 1.790 ;
        RECT  0.100 1.630 0.380 1.910 ;
        RECT  1.280 1.630 1.440 2.100 ;
        RECT  2.320 1.580 2.480 2.100 ;
        RECT  1.280 1.940 2.480 2.100 ;
        RECT  1.740 0.620 2.960 0.780 ;
        RECT  1.740 0.620 1.900 1.150 ;
        RECT  1.460 0.950 1.900 1.150 ;
        RECT  2.800 0.620 2.960 1.990 ;
        RECT  2.800 1.770 3.100 1.990 ;
        RECT  1.420 0.300 3.280 0.460 ;
        RECT  0.100 0.420 0.400 0.680 ;
        RECT  1.420 0.300 1.580 0.680 ;
        RECT  0.100 0.480 1.580 0.680 ;
        RECT  3.120 0.300 3.280 0.880 ;
        RECT  3.120 0.720 3.940 0.880 ;
        RECT  3.780 0.720 3.940 1.290 ;
        RECT  1.140 0.480 1.300 1.470 ;
        RECT  1.140 1.310 1.860 1.470 ;
        RECT  1.700 1.310 1.860 1.780 ;
        RECT  1.700 1.620 2.060 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO22B10M2HM

MACRO AO22B10M1HM
    CLASS CORE ;
    FOREIGN AO22B10M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.935  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.080 2.300 1.280 ;
        LAYER ME2 ;
        RECT  2.100 0.990 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.940 2.460 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.340 1.280 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.980 1.320 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.180 1.140 3.560 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.870 1.730 4.300 2.010 ;
        RECT  4.100 0.390 4.300 2.010 ;
        RECT  3.850 0.390 4.300 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.420 1.810 3.620 2.540 ;
        RECT  0.660 1.950 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.440 -0.140 3.640 0.650 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.630 1.440 1.790 ;
        RECT  0.100 1.630 0.380 1.910 ;
        RECT  1.280 1.630 1.440 2.100 ;
        RECT  2.320 1.580 2.480 2.100 ;
        RECT  1.280 1.940 2.480 2.100 ;
        RECT  1.740 0.620 2.960 0.780 ;
        RECT  1.740 0.620 1.900 1.150 ;
        RECT  1.460 0.950 1.900 1.150 ;
        RECT  2.800 0.620 2.960 2.010 ;
        RECT  2.800 1.810 3.100 2.010 ;
        RECT  1.420 0.300 3.280 0.460 ;
        RECT  0.100 0.420 0.400 0.680 ;
        RECT  1.420 0.300 1.580 0.680 ;
        RECT  0.100 0.480 1.580 0.680 ;
        RECT  3.120 0.300 3.280 0.970 ;
        RECT  3.120 0.810 3.940 0.970 ;
        RECT  3.780 0.810 3.940 1.290 ;
        RECT  1.140 0.480 1.300 1.470 ;
        RECT  1.140 1.310 1.860 1.470 ;
        RECT  1.700 1.310 1.860 1.780 ;
        RECT  1.700 1.620 2.060 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO22B10M1HM

MACRO AO22B10M0HM
    CLASS CORE ;
    FOREIGN AO22B10M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        ANTENNAGATEAREA 0.086  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.935  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.080 2.300 1.280 ;
        LAYER ME2 ;
        RECT  2.100 0.990 2.300 1.560 ;
        LAYER ME1 ;
        RECT  2.060 0.940 2.460 1.360 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.340 1.280 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.086  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 0.840 0.980 1.320 ;
        END
    END B2
    PIN NA2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.083  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.180 1.140 3.560 1.560 ;
        END
    END NA2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.870 1.730 4.300 2.010 ;
        RECT  4.100 0.390 4.300 2.010 ;
        RECT  3.850 0.390 4.300 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.420 1.810 3.620 2.540 ;
        RECT  0.660 1.950 0.940 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.440 -0.140 3.640 0.650 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.630 1.440 1.790 ;
        RECT  0.100 1.630 0.380 1.910 ;
        RECT  1.280 1.630 1.440 2.100 ;
        RECT  2.300 1.620 2.500 2.100 ;
        RECT  1.280 1.940 2.500 2.100 ;
        RECT  1.740 0.620 2.960 0.780 ;
        RECT  1.740 0.620 1.900 1.150 ;
        RECT  1.460 0.950 1.900 1.150 ;
        RECT  2.800 0.620 2.960 2.010 ;
        RECT  2.800 1.810 3.100 2.010 ;
        RECT  1.420 0.300 3.280 0.460 ;
        RECT  0.100 0.420 0.400 0.680 ;
        RECT  1.420 0.300 1.580 0.680 ;
        RECT  0.100 0.480 1.580 0.680 ;
        RECT  3.120 0.300 3.280 0.970 ;
        RECT  3.120 0.810 3.940 0.970 ;
        RECT  3.780 0.810 3.940 1.290 ;
        RECT  1.140 0.480 1.300 1.470 ;
        RECT  1.140 1.310 1.860 1.470 ;
        RECT  1.700 1.310 1.860 1.780 ;
        RECT  1.700 1.620 2.060 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO22B10M0HM

MACRO AO222M8HM
    CLASS CORE ;
    FOREIGN AO222M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        ANTENNAGATEAREA 0.286  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.620  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 0.840 3.500 1.040 ;
        LAYER ME2 ;
        RECT  3.300 0.680 3.500 1.320 ;
        LAYER ME1 ;
        RECT  3.040 0.820 3.680 1.070 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        ANTENNAGATEAREA 0.286  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.711  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 0.880 1.500 1.080 ;
        LAYER ME2 ;
        RECT  1.300 0.790 1.500 1.560 ;
        LAYER ME1 ;
        RECT  0.960 0.850 1.650 1.100 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.276  LAYER ME1  ;
        ANTENNAGATEAREA 0.276  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 0.850 5.900 1.050 ;
        LAYER ME2 ;
        RECT  5.700 0.690 5.900 1.380 ;
        LAYER ME1 ;
        RECT  5.600 0.820 6.240 1.070 ;
        END
    END C1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.260 2.020 1.420 ;
        RECT  1.860 0.900 2.020 1.420 ;
        RECT  0.500 0.840 0.700 1.420 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 1.230 4.100 1.390 ;
        RECT  3.940 0.890 4.100 1.390 ;
        RECT  2.500 0.810 2.740 1.390 ;
        END
    END B2
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.276  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.180 1.230 6.700 1.390 ;
        RECT  6.500 0.810 6.700 1.390 ;
        RECT  5.180 0.850 5.340 1.390 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.380 1.520 8.700 2.100 ;
        RECT  8.500 0.370 8.700 2.100 ;
        RECT  7.380 0.660 8.700 0.820 ;
        RECT  8.420 0.370 8.700 0.820 ;
        RECT  7.340 1.520 8.700 1.720 ;
        RECT  7.340 1.520 7.640 2.100 ;
        RECT  7.380 0.370 7.580 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.900 1.420 9.180 2.540 ;
        RECT  7.860 1.880 8.140 2.540 ;
        RECT  6.860 1.450 7.100 2.540 ;
        RECT  5.780 1.900 6.060 2.540 ;
        RECT  4.740 1.900 5.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.940 -0.140 9.140 0.710 ;
        RECT  7.860 -0.140 8.140 0.500 ;
        RECT  6.720 -0.140 7.000 0.320 ;
        RECT  4.900 -0.140 5.180 0.320 ;
        RECT  4.100 -0.140 4.380 0.320 ;
        RECT  2.180 -0.140 2.460 0.320 ;
        RECT  0.340 -0.140 0.540 0.630 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.440 0.340 2.100 ;
        RECT  1.140 1.900 1.420 2.100 ;
        RECT  2.180 1.900 2.460 2.100 ;
        RECT  3.220 1.900 3.510 2.100 ;
        RECT  4.220 1.900 4.540 2.100 ;
        RECT  0.140 1.940 4.540 2.100 ;
        RECT  2.620 1.560 6.580 1.720 ;
        RECT  5.260 1.560 5.540 1.980 ;
        RECT  6.300 1.560 6.580 1.980 ;
        RECT  1.100 0.480 7.220 0.640 ;
        RECT  7.060 0.480 7.220 1.240 ;
        RECT  7.060 1.040 8.300 1.240 ;
        RECT  2.180 0.480 2.340 1.740 ;
        RECT  0.590 1.580 2.340 1.740 ;
        RECT  0.590 1.580 0.950 1.780 ;
        RECT  1.610 1.580 1.970 1.780 ;
        LAYER VTPH ;
        RECT  1.500 1.050 4.860 2.400 ;
        RECT  0.000 1.080 4.860 2.400 ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.050 ;
        RECT  0.000 0.000 1.500 1.080 ;
        RECT  4.860 0.000 9.600 1.140 ;
    END
END AO222M8HM

MACRO AO222M4HM
    CLASS CORE ;
    FOREIGN AO222M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.380 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.320 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 0.840 1.900 1.250 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.060 0.840 2.300 1.300 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.080 0.840 3.500 1.320 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 1.040 3.900 1.560 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.300 1.480 5.100 1.680 ;
        RECT  4.900 0.680 5.100 1.680 ;
        RECT  4.460 0.680 5.100 0.880 ;
        RECT  4.460 0.360 4.660 0.880 ;
        RECT  4.300 1.480 4.580 2.060 ;
        RECT  4.300 0.360 4.660 0.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.820 1.840 5.100 2.540 ;
        RECT  3.780 1.800 4.060 2.540 ;
        RECT  2.740 1.900 3.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.820 -0.140 5.100 0.520 ;
        RECT  3.740 -0.140 4.020 0.320 ;
        RECT  2.220 -0.140 2.500 0.320 ;
        RECT  0.140 -0.140 0.340 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.540 0.380 2.100 ;
        RECT  1.140 1.540 1.420 2.100 ;
        RECT  2.180 1.900 2.460 2.100 ;
        RECT  0.100 1.940 2.460 2.100 ;
        RECT  1.620 1.580 3.400 1.740 ;
        RECT  1.620 1.580 1.970 1.780 ;
        RECT  3.220 1.580 3.400 1.970 ;
        RECT  3.220 1.810 3.600 1.970 ;
        RECT  0.540 0.480 3.970 0.640 ;
        RECT  3.800 0.480 3.970 0.880 ;
        RECT  3.800 0.720 4.260 0.880 ;
        RECT  4.100 0.720 4.260 1.320 ;
        RECT  4.100 1.040 4.720 1.320 ;
        RECT  0.540 0.480 0.700 1.760 ;
        RECT  0.540 1.600 0.940 1.760 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END AO222M4HM

MACRO AO222M2HM
    CLASS CORE ;
    FOREIGN AO222M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.120 1.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.900 1.980 1.320 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 0.840 2.740 1.250 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.160 0.840 3.500 1.320 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 1.040 3.900 1.590 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.410 4.700 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.840 -0.140 4.120 0.320 ;
        RECT  2.380 -0.140 2.660 0.320 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.790 0.340 2.100 ;
        RECT  1.260 1.790 1.460 2.100 ;
        RECT  2.280 1.900 2.670 2.100 ;
        RECT  0.140 1.940 2.670 2.100 ;
        RECT  1.690 1.580 3.460 1.740 ;
        RECT  1.690 1.580 2.110 1.780 ;
        RECT  3.300 1.580 3.460 2.060 ;
        RECT  3.300 1.900 3.700 2.060 ;
        RECT  0.580 0.480 4.300 0.640 ;
        RECT  4.140 0.480 4.300 1.360 ;
        RECT  0.580 0.480 0.740 1.780 ;
        RECT  0.580 1.620 1.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO222M2HM

MACRO AO222M1HM
    CLASS CORE ;
    FOREIGN AO222M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.120 1.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.640 0.900 1.980 1.320 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 0.840 2.740 1.300 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.160 0.840 3.500 1.320 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 1.040 3.900 1.590 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.410 4.700 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.840 -0.140 4.120 0.320 ;
        RECT  2.380 -0.140 2.660 0.320 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.790 0.340 2.100 ;
        RECT  1.260 1.790 1.460 2.100 ;
        RECT  2.280 1.900 2.670 2.100 ;
        RECT  0.140 1.940 2.670 2.100 ;
        RECT  1.690 1.580 3.460 1.740 ;
        RECT  1.690 1.580 2.110 1.780 ;
        RECT  3.300 1.580 3.460 2.060 ;
        RECT  3.300 1.900 3.700 2.060 ;
        RECT  0.580 0.480 4.300 0.640 ;
        RECT  4.140 0.480 4.300 1.360 ;
        RECT  0.580 0.480 0.740 1.780 ;
        RECT  0.580 1.620 1.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO222M1HM

MACRO AO222M0HM
    CLASS CORE ;
    FOREIGN AO222M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.220 1.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.560 0.900 1.980 1.280 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.220 0.840 2.700 1.250 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.160 0.840 3.500 1.320 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.096  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.660 1.040 3.900 1.590 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.480 0.410 4.700 2.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  3.900 1.900 4.180 2.540 ;
        RECT  2.860 1.900 3.140 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  3.840 -0.140 4.120 0.320 ;
        RECT  2.380 -0.140 2.660 0.320 ;
        RECT  0.140 -0.140 0.340 0.680 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 1.790 0.340 2.100 ;
        RECT  1.260 1.790 1.460 2.100 ;
        RECT  2.280 1.900 2.670 2.100 ;
        RECT  0.140 1.940 2.670 2.100 ;
        RECT  1.690 1.580 3.460 1.740 ;
        RECT  1.690 1.580 2.110 1.780 ;
        RECT  3.300 1.580 3.460 2.060 ;
        RECT  3.300 1.900 3.700 2.060 ;
        RECT  0.580 0.480 4.300 0.640 ;
        RECT  4.140 0.480 4.300 1.360 ;
        RECT  0.580 0.480 0.740 1.780 ;
        RECT  0.580 1.620 1.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO222M0HM

MACRO AO221M8HM
    CLASS CORE ;
    FOREIGN AO221M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.244  LAYER ME1  ;
        ANTENNAGATEAREA 0.244  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.049  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.500 1.080 0.700 1.280 ;
        LAYER ME2 ;
        RECT  0.500 0.940 0.700 1.600 ;
        LAYER ME1 ;
        RECT  0.440 1.040 1.100 1.340 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME2  ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.529  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 0.860 2.700 1.060 ;
        LAYER ME2 ;
        RECT  2.500 0.720 2.700 1.380 ;
        LAYER ME1 ;
        RECT  2.150 0.850 2.760 1.080 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        ANTENNAGATEAREA 0.286  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.730  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.900 0.860 5.100 1.060 ;
        LAYER ME2 ;
        RECT  4.900 0.720 5.100 1.560 ;
        LAYER ME1 ;
        RECT  4.440 0.850 5.160 1.080 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.240 5.660 1.400 ;
        RECT  5.500 0.850 5.660 1.400 ;
        RECT  4.100 0.900 4.260 1.400 ;
        RECT  3.640 0.900 4.260 1.110 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.286  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 1.240 3.100 1.400 ;
        RECT  2.940 0.930 3.100 1.400 ;
        RECT  1.540 0.840 1.960 1.400 ;
        END
    END B1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.860 0.370 8.060 2.100 ;
        RECT  6.780 1.520 8.060 1.720 ;
        RECT  7.700 0.660 8.060 1.720 ;
        RECT  6.820 0.660 8.060 0.840 ;
        RECT  6.780 1.520 7.020 2.100 ;
        RECT  6.820 0.370 7.020 0.840 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.800 2.540 ;
        RECT  8.380 1.460 8.580 2.540 ;
        RECT  7.300 1.880 7.580 2.540 ;
        RECT  6.300 1.460 6.500 2.540 ;
        RECT  0.620 1.880 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.800 0.140 ;
        RECT  8.380 -0.140 8.580 0.650 ;
        RECT  7.300 -0.140 7.580 0.500 ;
        RECT  6.260 -0.140 6.460 0.690 ;
        RECT  4.740 -0.140 5.020 0.340 ;
        RECT  2.180 -0.140 2.460 0.320 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.260 1.400 3.520 1.720 ;
        RECT  0.140 1.560 3.520 1.720 ;
        RECT  0.140 1.560 0.340 2.100 ;
        RECT  1.180 1.560 1.380 2.100 ;
        RECT  1.620 1.880 5.580 2.040 ;
        RECT  2.980 0.370 4.580 0.530 ;
        RECT  1.060 0.480 3.140 0.640 ;
        RECT  0.140 0.300 0.340 0.820 ;
        RECT  5.620 0.350 6.020 0.690 ;
        RECT  4.420 0.530 6.020 0.690 ;
        RECT  1.060 0.480 1.220 0.820 ;
        RECT  0.140 0.660 1.220 0.820 ;
        RECT  5.820 1.040 7.500 1.240 ;
        RECT  3.680 1.400 3.940 1.720 ;
        RECT  3.680 1.560 6.020 1.720 ;
        RECT  5.820 0.350 6.020 2.100 ;
        LAYER VTPH ;
        RECT  0.440 1.100 6.220 2.400 ;
        RECT  0.000 1.140 8.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.800 1.100 ;
        RECT  0.000 0.000 0.440 1.140 ;
        RECT  6.220 0.000 8.800 1.140 ;
    END
END AO221M8HM

MACRO AO221M4HM
    CLASS CORE ;
    FOREIGN AO221M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.900 1.560 1.340 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 0.840 0.700 1.300 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 1.060 3.100 1.560 ;
        RECT  2.600 1.060 3.100 1.260 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.900 2.360 1.300 ;
        END
    END B2
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 1.020 3.500 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.900 1.540 4.700 1.740 ;
        RECT  4.500 0.680 4.700 1.740 ;
        RECT  4.020 0.680 4.700 0.880 ;
        RECT  4.020 0.340 4.220 0.880 ;
        RECT  3.900 1.540 4.190 2.100 ;
        RECT  3.900 0.340 4.220 0.540 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.420 1.900 4.700 2.540 ;
        RECT  3.380 1.900 3.660 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.420 -0.140 4.700 0.520 ;
        RECT  3.340 -0.140 3.620 0.320 ;
        RECT  1.900 -0.140 2.180 0.320 ;
        RECT  0.340 -0.140 0.540 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 1.580 2.660 1.740 ;
        RECT  0.100 1.540 0.380 2.100 ;
        RECT  1.200 1.580 1.360 2.100 ;
        RECT  0.100 1.940 1.360 2.100 ;
        RECT  1.780 1.900 3.180 2.060 ;
        RECT  0.860 0.540 3.560 0.700 ;
        RECT  3.400 0.700 3.820 0.860 ;
        RECT  3.660 0.700 3.820 1.320 ;
        RECT  3.660 1.040 4.320 1.320 ;
        RECT  0.860 0.540 1.020 1.780 ;
        RECT  0.580 1.620 1.020 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AO221M4HM

MACRO AO221M2HM
    CLASS CORE ;
    FOREIGN AO221M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.840 3.500 1.340 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.900 1.560 1.390 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 0.840 0.700 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.600 0.840 3.100 1.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.900 2.360 1.400 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.410 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.500 1.500 3.780 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.460 -0.140 3.740 0.320 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.340 -0.140 0.540 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 1.560 2.780 1.720 ;
        RECT  0.100 1.520 0.380 2.040 ;
        RECT  1.200 1.560 1.360 2.040 ;
        RECT  0.100 1.880 1.360 2.040 ;
        RECT  1.900 1.880 3.300 2.040 ;
        RECT  0.860 0.510 3.900 0.670 ;
        RECT  3.740 0.510 3.900 1.340 ;
        RECT  0.860 0.510 1.020 1.720 ;
        RECT  0.580 1.560 1.020 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO221M2HM

MACRO AO221M1HM
    CLASS CORE ;
    FOREIGN AO221M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.840 3.500 1.340 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.900 1.560 1.390 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 0.840 0.700 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.600 0.840 3.100 1.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.900 2.360 1.400 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.410 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.540 1.760 3.740 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.460 -0.140 3.740 0.320 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.340 -0.140 0.540 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 1.560 2.780 1.720 ;
        RECT  0.100 1.520 0.380 2.040 ;
        RECT  1.200 1.560 1.360 2.040 ;
        RECT  0.100 1.880 1.360 2.040 ;
        RECT  1.900 1.880 3.300 2.040 ;
        RECT  0.860 0.510 3.900 0.670 ;
        RECT  3.740 0.510 3.900 1.340 ;
        RECT  0.860 0.510 1.020 1.720 ;
        RECT  0.580 1.560 1.020 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO221M1HM

MACRO AO221M0HM
    CLASS CORE ;
    FOREIGN AO221M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.260 0.840 3.500 1.340 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.180 0.900 1.560 1.390 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 0.840 0.700 1.360 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.600 0.840 3.100 1.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.040 0.900 2.360 1.400 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.080 0.410 4.300 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.500 1.700 3.780 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.460 -0.140 3.740 0.320 ;
        RECT  2.020 -0.140 2.300 0.320 ;
        RECT  0.340 -0.140 0.540 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 1.560 2.780 1.720 ;
        RECT  0.100 1.520 0.380 2.040 ;
        RECT  1.200 1.560 1.360 2.040 ;
        RECT  0.100 1.880 1.360 2.040 ;
        RECT  1.900 1.880 3.300 2.040 ;
        RECT  0.860 0.510 3.900 0.670 ;
        RECT  3.740 0.510 3.900 1.340 ;
        RECT  0.860 0.510 1.020 1.720 ;
        RECT  0.580 1.560 1.020 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.400 1.140 ;
    END
END AO221M0HM

MACRO AO21M8HM
    CLASS CORE ;
    FOREIGN AO21M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.250  LAYER ME1  ;
        ANTENNAGATEAREA 0.250  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.833  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.040 3.500 1.240 ;
        LAYER ME2 ;
        RECT  3.300 0.900 3.500 1.560 ;
        LAYER ME1 ;
        RECT  3.080 1.000 3.680 1.280 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.282  LAYER ME1  ;
        ANTENNAGATEAREA 0.282  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.826  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.080 1.500 1.280 ;
        LAYER ME2 ;
        RECT  1.300 1.020 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.200 1.020 1.870 1.300 ;
        RECT  1.300 1.020 1.500 1.340 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.284  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.020 1.040 1.300 ;
        RECT  0.100 1.020 0.300 1.560 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.340 0.660 5.620 2.100 ;
        RECT  5.380 0.390 5.620 2.100 ;
        RECT  4.300 1.540 5.620 1.740 ;
        RECT  5.290 0.660 5.620 1.740 ;
        RECT  4.340 0.660 5.620 0.860 ;
        RECT  4.300 1.540 4.600 2.100 ;
        RECT  4.340 0.390 4.540 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.400 2.540 ;
        RECT  5.900 1.480 6.100 2.540 ;
        RECT  4.820 1.900 5.100 2.540 ;
        RECT  3.780 1.900 4.060 2.540 ;
        RECT  2.700 2.080 2.980 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.400 0.140 ;
        RECT  5.900 -0.140 6.100 0.690 ;
        RECT  4.820 -0.140 5.100 0.500 ;
        RECT  3.780 -0.140 4.060 0.500 ;
        RECT  2.740 -0.140 3.020 0.500 ;
        RECT  0.620 -0.140 0.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.200 0.320 2.580 0.480 ;
        RECT  2.160 0.320 2.580 0.500 ;
        RECT  0.140 0.370 0.340 0.820 ;
        RECT  1.200 0.320 1.360 0.820 ;
        RECT  0.140 0.660 1.360 0.820 ;
        RECT  0.100 1.810 0.380 2.050 ;
        RECT  2.340 1.760 3.580 1.920 ;
        RECT  0.100 1.890 2.500 2.050 ;
        RECT  1.660 0.640 2.020 0.820 ;
        RECT  3.300 0.310 3.500 0.820 ;
        RECT  1.660 0.660 4.140 0.820 ;
        RECT  3.980 1.040 5.120 1.250 ;
        RECT  2.020 1.440 4.140 1.600 ;
        RECT  3.980 0.660 4.140 1.600 ;
        RECT  0.580 1.570 2.180 1.730 ;
        LAYER VTPH ;
        RECT  0.000 1.140 1.480 2.400 ;
        RECT  2.160 1.140 6.400 2.400 ;
        RECT  0.000 1.160 6.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.400 1.140 ;
        RECT  1.480 0.000 2.160 1.160 ;
    END
END AO21M8HM

MACRO AO21M4HM
    CLASS CORE ;
    FOREIGN AO21M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.127  LAYER ME1  ;
        ANTENNAGATEAREA 0.127  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.516  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.060 1.500 1.260 ;
        LAYER ME2 ;
        RECT  1.300 0.870 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.260 0.980 1.760 1.340 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.620 1.100 1.300 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.145  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.300 0.840 0.700 1.310 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.300 1.520 3.100 1.720 ;
        RECT  2.900 0.660 3.100 1.720 ;
        RECT  2.360 0.660 3.100 0.820 ;
        RECT  2.300 1.520 2.600 2.100 ;
        RECT  2.360 0.410 2.580 0.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 1.900 3.100 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.500 ;
        RECT  1.780 -0.140 2.060 0.500 ;
        RECT  0.260 -0.140 0.460 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.220 1.530 0.500 2.060 ;
        RECT  0.220 1.900 1.620 2.060 ;
        RECT  1.260 0.400 1.460 0.820 ;
        RECT  1.260 0.660 2.140 0.820 ;
        RECT  1.940 1.040 2.720 1.320 ;
        RECT  1.940 0.660 2.140 1.740 ;
        RECT  0.690 1.580 2.140 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO21M4HM

MACRO AO21M2HM
    CLASS CORE ;
    FOREIGN AO21M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.560 1.040 1.960 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.080 1.280 1.280 ;
        RECT  0.900 0.840 1.160 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.450 0.840 0.740 1.250 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.480 0.410 2.700 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.520 ;
        RECT  0.380 -0.140 0.580 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 1.690 0.580 2.100 ;
        RECT  1.300 1.900 1.690 2.100 ;
        RECT  0.380 1.940 1.690 2.100 ;
        RECT  1.320 0.350 1.520 0.840 ;
        RECT  1.320 0.680 2.320 0.840 ;
        RECT  2.120 0.680 2.320 1.740 ;
        RECT  0.860 1.580 2.320 1.740 ;
        RECT  0.860 1.580 1.140 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AO21M2HM

MACRO AO21M1HM
    CLASS CORE ;
    FOREIGN AO21M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.560 1.040 1.960 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.080 1.280 1.280 ;
        RECT  0.900 0.440 1.100 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.740 1.250 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.480 0.350 2.700 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.520 ;
        RECT  0.380 -0.140 0.580 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 1.690 0.580 2.100 ;
        RECT  1.300 1.900 1.690 2.100 ;
        RECT  0.380 1.940 1.690 2.100 ;
        RECT  1.320 0.350 1.520 0.880 ;
        RECT  1.320 0.680 2.320 0.880 ;
        RECT  2.120 0.680 2.320 1.740 ;
        RECT  0.830 1.580 2.320 1.740 ;
        RECT  0.830 1.580 1.140 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AO21M1HM

MACRO AO21M0HM
    CLASS CORE ;
    FOREIGN AO21M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.106  LAYER ME1  ;
        ANTENNAGATEAREA 0.106  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.841  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.140 1.900 1.340 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.560 1.040 1.960 1.420 ;
        END
    END B
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.080 1.280 1.280 ;
        RECT  0.900 0.440 1.100 1.280 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.121  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.340 0.840 0.740 1.250 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.480 0.300 2.700 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.900 1.900 2.180 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.900 -0.140 2.180 0.520 ;
        RECT  0.380 -0.140 0.580 0.620 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.380 1.690 0.580 2.100 ;
        RECT  1.300 1.900 1.690 2.100 ;
        RECT  0.380 1.940 1.690 2.100 ;
        RECT  1.320 0.350 1.520 0.880 ;
        RECT  1.320 0.680 2.320 0.880 ;
        RECT  2.120 0.680 2.320 1.740 ;
        RECT  0.830 1.580 2.320 1.740 ;
        RECT  0.830 1.580 1.140 1.780 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AO21M0HM

MACRO AO211M8HM
    CLASS CORE ;
    FOREIGN AO211M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME2  ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 1.807  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.060 1.500 1.260 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.400 ;
        LAYER ME1 ;
        RECT  1.080 1.040 1.720 1.280 ;
        END
    END C
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.276  LAYER ME1  ;
        ANTENNAGATEAREA 0.276  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.130 3.500 1.330 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.400 ;
        LAYER ME1 ;
        RECT  3.040 1.120 3.680 1.370 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.276  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.980 0.800 4.140 1.320 ;
        RECT  2.500 0.800 4.140 0.960 ;
        RECT  2.500 0.800 2.740 1.400 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.253  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 2.180 1.600 ;
        RECT  1.980 1.000 2.180 1.600 ;
        RECT  0.500 1.000 0.740 1.600 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.500 0.660 6.700 1.740 ;
        RECT  6.300 1.540 6.580 2.100 ;
        RECT  6.340 0.390 6.540 0.880 ;
        RECT  5.300 0.660 6.700 0.880 ;
        RECT  5.260 1.540 6.700 1.720 ;
        RECT  5.260 1.540 5.540 2.100 ;
        RECT  5.300 0.390 5.500 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.860 1.480 7.060 2.540 ;
        RECT  5.780 1.900 6.060 2.540 ;
        RECT  4.800 1.450 5.000 2.540 ;
        RECT  1.220 2.080 1.500 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.860 -0.140 7.060 0.660 ;
        RECT  5.780 -0.140 6.060 0.500 ;
        RECT  4.800 -0.140 5.000 0.670 ;
        RECT  4.100 -0.140 4.380 0.320 ;
        RECT  2.340 -0.140 2.620 0.320 ;
        RECT  1.260 -0.140 1.540 0.500 ;
        RECT  0.260 -0.140 0.460 0.570 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.300 1.760 2.470 1.920 ;
        RECT  2.310 1.900 4.580 2.060 ;
        RECT  1.780 0.300 2.060 0.640 ;
        RECT  1.780 0.480 4.640 0.640 ;
        RECT  0.740 0.300 1.020 0.840 ;
        RECT  1.780 0.300 2.000 0.840 ;
        RECT  0.740 0.660 2.000 0.840 ;
        RECT  4.480 1.080 6.340 1.280 ;
        RECT  4.480 0.480 4.640 1.740 ;
        RECT  2.660 1.580 4.640 1.740 ;
        LAYER VTPH ;
        RECT  0.000 1.050 4.500 2.400 ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.050 ;
        RECT  4.500 0.000 7.200 1.140 ;
    END
END AO211M8HM

MACRO AO211M4HM
    CLASS CORE ;
    FOREIGN AO211M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.310 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.138  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.310 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.950 1.500 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.990 2.040 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.540 3.500 1.740 ;
        RECT  3.300 0.660 3.500 1.740 ;
        RECT  2.700 0.660 3.500 0.860 ;
        RECT  2.660 1.540 2.940 2.100 ;
        RECT  2.700 0.390 2.900 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.180 1.900 3.460 2.540 ;
        RECT  2.060 1.880 2.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.180 -0.140 3.460 0.500 ;
        RECT  2.100 -0.140 2.380 0.320 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.540 0.380 2.060 ;
        RECT  0.100 1.900 1.460 2.060 ;
        RECT  0.140 0.340 0.340 0.640 ;
        RECT  1.540 0.300 1.820 0.640 ;
        RECT  0.140 0.480 2.540 0.640 ;
        RECT  2.380 0.480 2.540 1.280 ;
        RECT  2.380 1.080 3.120 1.280 ;
        RECT  0.540 0.480 0.700 1.720 ;
        RECT  0.540 1.560 0.940 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AO211M4HM

MACRO AO211M2HM
    CLASS CORE ;
    FOREIGN AO211M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.310 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.310 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.950 1.500 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.990 2.040 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.540 3.100 2.100 ;
        RECT  2.900 0.660 3.100 2.100 ;
        RECT  2.700 0.390 2.900 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.060 1.880 2.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.100 -0.140 2.380 0.320 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.540 0.380 2.060 ;
        RECT  0.100 1.900 1.460 2.060 ;
        RECT  0.140 0.340 0.340 0.640 ;
        RECT  1.540 0.300 1.820 0.640 ;
        RECT  0.140 0.480 2.540 0.640 ;
        RECT  2.380 0.480 2.540 1.360 ;
        RECT  0.540 0.480 0.700 1.720 ;
        RECT  0.540 1.560 0.940 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO211M2HM

MACRO AO211M1HM
    CLASS CORE ;
    FOREIGN AO211M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.310 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.310 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.950 1.500 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.990 2.040 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.540 3.100 1.740 ;
        RECT  2.900 0.660 3.100 1.740 ;
        RECT  2.700 0.390 2.900 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.060 1.880 2.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.100 -0.140 2.380 0.320 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.540 0.380 2.060 ;
        RECT  0.100 1.900 1.460 2.060 ;
        RECT  0.140 0.340 0.340 0.640 ;
        RECT  1.540 0.300 1.820 0.640 ;
        RECT  0.140 0.480 2.540 0.640 ;
        RECT  2.380 0.480 2.540 1.360 ;
        RECT  0.540 0.480 0.700 1.720 ;
        RECT  0.540 1.560 0.940 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO211M1HM

MACRO AO211M0HM
    CLASS CORE ;
    FOREIGN AO211M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.380 1.310 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.400 ;
        END
    END A2
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.950 1.500 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 0.990 2.040 1.560 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.660 1.680 3.100 1.880 ;
        RECT  2.900 0.660 3.100 1.880 ;
        RECT  2.700 0.390 2.900 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.060 1.880 2.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.100 -0.140 2.380 0.320 ;
        RECT  0.980 -0.140 1.260 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 1.540 0.380 2.060 ;
        RECT  0.100 1.900 1.460 2.060 ;
        RECT  0.140 0.340 0.340 0.640 ;
        RECT  1.540 0.300 1.820 0.640 ;
        RECT  0.140 0.480 2.540 0.640 ;
        RECT  2.380 0.480 2.540 1.360 ;
        RECT  0.540 0.480 0.700 1.720 ;
        RECT  0.540 1.560 0.940 1.720 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AO211M0HM

MACRO ANTHM
    CLASS CORE ;
    FOREIGN ANTHM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.372  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.430 0.540 0.630 ;
        RECT  0.100 0.430 0.300 1.160 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 0.800 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 0.800 0.140 ;
        END
    END VSS
    OBS
        LAYER VTPH ;
        RECT  0.000 1.140 0.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 0.800 1.140 ;
    END
END ANTHM

MACRO AN4M8HM
    CLASS CORE ;
    FOREIGN AN4M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME2  ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 2.145  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  3.300 1.010 3.500 1.210 ;
        LAYER ME2 ;
        RECT  3.300 0.840 3.500 1.400 ;
        LAYER ME1 ;
        RECT  3.160 0.990 3.880 1.240 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        ANTENNAGATEAREA 0.235  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.968  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.140 1.500 1.340 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.400 ;
        LAYER ME1 ;
        RECT  1.000 1.120 1.640 1.370 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.680 1.430 4.300 1.590 ;
        RECT  4.100 1.050 4.300 1.590 ;
        RECT  2.680 1.090 2.880 1.590 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.900 0.800 2.100 1.370 ;
        RECT  0.500 0.800 2.100 0.960 ;
        RECT  0.500 0.800 0.700 1.410 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.300 1.540 6.700 2.100 ;
        RECT  6.500 0.390 6.700 2.100 ;
        RECT  5.300 0.660 6.700 0.860 ;
        RECT  6.360 0.390 6.700 0.860 ;
        RECT  5.260 1.540 6.700 1.740 ;
        RECT  5.260 1.540 5.550 2.100 ;
        RECT  5.300 0.390 5.500 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.860 1.480 7.060 2.540 ;
        RECT  5.780 1.900 6.060 2.540 ;
        RECT  4.600 2.080 4.880 2.540 ;
        RECT  3.380 2.080 3.660 2.540 ;
        RECT  2.260 2.080 2.540 2.540 ;
        RECT  1.180 1.900 1.460 2.540 ;
        RECT  0.180 1.770 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.860 -0.140 7.060 0.650 ;
        RECT  5.780 -0.140 6.060 0.500 ;
        RECT  4.740 -0.140 5.020 0.500 ;
        RECT  1.140 -0.140 1.420 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.620 0.300 4.540 0.460 ;
        RECT  4.260 0.300 4.540 0.500 ;
        RECT  2.620 0.300 2.820 0.640 ;
        RECT  0.220 0.480 2.820 0.640 ;
        RECT  3.330 0.620 3.660 0.820 ;
        RECT  3.330 0.660 5.100 0.820 ;
        RECT  4.900 1.080 6.300 1.280 ;
        RECT  0.720 1.580 1.800 1.740 ;
        RECT  1.640 1.580 1.800 1.920 ;
        RECT  4.900 0.660 5.100 1.920 ;
        RECT  1.640 1.760 5.100 1.920 ;
        RECT  0.720 1.580 0.880 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END AN4M8HM

MACRO AN4M6HM
    CLASS CORE ;
    FOREIGN AN4M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER ME1  ;
        ANTENNAGATEAREA 0.200  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.425  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.500 1.100 1.700 ;
        LAYER ME2 ;
        RECT  0.900 1.240 1.100 1.800 ;
        LAYER ME1 ;
        RECT  0.840 1.440 1.820 1.600 ;
        RECT  0.840 1.440 1.100 1.780 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER ME1  ;
        ANTENNAGATEAREA 0.200  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.086  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.100 1.000 2.300 1.200 ;
        LAYER ME2 ;
        RECT  2.100 0.830 2.300 1.560 ;
        LAYER ME1 ;
        RECT  1.240 0.960 2.960 1.200 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 0.620 3.500 1.240 ;
        RECT  0.820 0.620 3.500 0.780 ;
        RECT  0.820 0.620 0.980 1.230 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.980 1.440 3.900 1.600 ;
        RECT  3.700 1.040 3.900 1.600 ;
        RECT  1.460 1.760 2.140 1.920 ;
        RECT  1.980 1.440 2.140 1.920 ;
        RECT  0.340 1.940 1.620 2.100 ;
        RECT  1.460 1.760 1.620 2.100 ;
        RECT  0.340 0.850 0.500 2.100 ;
        END
    END D
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.620 1.540 5.900 2.100 ;
        RECT  5.700 0.390 5.900 2.100 ;
        RECT  4.620 0.660 5.900 0.860 ;
        RECT  5.680 0.390 5.900 0.860 ;
        RECT  4.580 1.540 5.900 1.740 ;
        RECT  4.580 1.540 4.860 2.100 ;
        RECT  4.620 0.390 4.820 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.100 1.900 5.380 2.540 ;
        RECT  4.020 2.080 4.300 2.540 ;
        RECT  2.900 2.080 3.180 2.540 ;
        RECT  1.780 2.080 2.060 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.100 -0.140 5.380 0.500 ;
        RECT  3.990 -0.140 4.270 0.320 ;
        RECT  0.140 -0.140 0.340 0.640 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.920 0.300 3.820 0.460 ;
        RECT  3.660 0.300 3.820 0.680 ;
        RECT  3.660 0.520 4.420 0.680 ;
        RECT  4.220 1.080 5.400 1.280 ;
        RECT  4.220 0.520 4.420 1.920 ;
        RECT  2.300 1.760 4.420 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END AN4M6HM

MACRO AN4M4HM
    CLASS CORE ;
    FOREIGN AN4M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        ANTENNAGATEAREA 0.118  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.449  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.130 1.900 1.330 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.700 1.040 2.100 1.420 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.118  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.700 1.540 3.500 1.740 ;
        RECT  3.300 0.660 3.500 1.740 ;
        RECT  2.740 0.660 3.500 0.860 ;
        RECT  2.700 1.540 2.980 2.100 ;
        RECT  2.740 0.390 2.940 0.860 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  3.220 -0.140 3.500 0.500 ;
        RECT  2.100 -0.140 2.380 0.500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.770 0.340 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.180 0.440 1.940 0.640 ;
        RECT  1.740 0.440 1.940 0.860 ;
        RECT  1.740 0.660 2.540 0.860 ;
        RECT  2.340 1.040 3.140 1.320 ;
        RECT  2.340 0.660 2.540 1.740 ;
        RECT  0.660 1.580 2.540 1.740 ;
        RECT  0.660 1.580 0.860 2.040 ;
        RECT  1.700 1.580 1.900 2.040 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AN4M4HM

MACRO AN4M2HM
    CLASS CORE ;
    FOREIGN AN4M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        ANTENNAGATEAREA 0.080  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.045  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.130 1.900 1.330 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.700 1.040 2.100 1.420 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.460 3.100 2.100 ;
        RECT  2.900 0.400 3.100 2.100 ;
        RECT  2.700 0.400 3.100 0.600 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.100 -0.140 2.380 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 0.440 1.940 0.640 ;
        RECT  1.740 0.440 1.940 0.860 ;
        RECT  1.740 0.660 2.540 0.860 ;
        RECT  2.340 0.660 2.540 1.740 ;
        RECT  0.620 1.580 2.540 1.740 ;
        RECT  0.620 1.580 0.900 2.100 ;
        RECT  1.660 1.580 1.940 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AN4M2HM

MACRO AN4M1HM
    CLASS CORE ;
    FOREIGN AN4M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        ANTENNAGATEAREA 0.080  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.045  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.130 1.900 1.330 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.700 1.040 2.100 1.420 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.700 1.880 3.100 2.080 ;
        RECT  2.900 0.380 3.100 2.080 ;
        RECT  2.700 0.380 3.100 0.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.100 -0.140 2.380 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 0.440 1.940 0.640 ;
        RECT  1.740 0.440 1.940 0.860 ;
        RECT  1.740 0.660 2.540 0.860 ;
        RECT  2.340 0.660 2.540 1.740 ;
        RECT  0.620 1.580 2.540 1.740 ;
        RECT  0.620 1.580 0.900 2.100 ;
        RECT  1.660 1.580 1.940 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AN4M1HM

MACRO AN4M16HM
    CLASS CORE ;
    FOREIGN AN4M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.130 1.100 1.330 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.520 1.080 1.520 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.080 1.080 3.080 1.400 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  10.020 1.540 10.300 2.100 ;
        RECT  6.940 0.680 10.260 0.880 ;
        RECT  10.060 0.410 10.260 0.880 ;
        RECT  6.900 1.540 10.300 1.740 ;
        RECT  8.980 1.540 9.260 2.100 ;
        RECT  9.020 0.410 9.220 0.880 ;
        RECT  8.500 0.680 8.750 1.740 ;
        RECT  7.940 1.540 8.220 2.100 ;
        RECT  7.980 0.410 8.180 0.880 ;
        RECT  6.900 1.540 7.180 2.100 ;
        RECT  6.940 0.410 7.140 0.880 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.130 4.300 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.400 ;
        LAYER ME1 ;
        RECT  3.640 1.080 4.640 1.400 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.130 5.900 1.330 ;
        LAYER ME2 ;
        RECT  5.700 0.840 5.900 1.400 ;
        LAYER ME1 ;
        RECT  5.200 1.080 6.200 1.400 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 11.200 2.540 ;
        RECT  10.540 1.540 10.820 2.540 ;
        RECT  9.500 1.900 9.780 2.540 ;
        RECT  8.460 1.900 8.740 2.540 ;
        RECT  7.420 1.900 7.700 2.540 ;
        RECT  6.360 1.900 6.640 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.710 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 11.200 0.140 ;
        RECT  10.540 -0.140 10.820 0.520 ;
        RECT  9.500 -0.140 9.780 0.520 ;
        RECT  8.460 -0.140 8.740 0.520 ;
        RECT  7.420 -0.140 7.700 0.520 ;
        RECT  6.400 -0.140 6.600 0.710 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.300 2.980 0.460 ;
        RECT  0.620 0.300 0.900 0.520 ;
        RECT  1.660 0.300 1.940 0.520 ;
        RECT  2.700 0.300 2.980 0.520 ;
        RECT  3.260 0.300 3.460 0.880 ;
        RECT  2.170 0.680 4.540 0.880 ;
        RECT  3.740 0.300 5.000 0.460 ;
        RECT  3.740 0.300 4.020 0.520 ;
        RECT  4.780 0.300 5.000 0.880 ;
        RECT  5.860 0.430 6.060 0.880 ;
        RECT  4.780 0.680 6.060 0.880 ;
        RECT  0.140 0.430 0.340 0.880 ;
        RECT  0.140 0.680 1.900 0.880 ;
        RECT  6.540 1.080 8.300 1.280 ;
        RECT  6.540 1.080 6.740 1.740 ;
        RECT  0.660 1.580 6.740 1.740 ;
        RECT  0.660 1.580 0.860 1.990 ;
        RECT  1.700 0.680 1.900 1.990 ;
        RECT  2.740 1.580 2.940 1.990 ;
        RECT  3.780 1.580 3.980 1.990 ;
        RECT  4.820 1.580 5.020 1.990 ;
        RECT  5.860 1.580 6.060 1.990 ;
        RECT  9.040 1.080 10.480 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.470 2.400 ;
        RECT  6.250 1.140 11.200 2.400 ;
        RECT  0.000 1.290 11.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 11.200 1.140 ;
        RECT  0.470 0.000 6.250 1.290 ;
    END
END AN4M16HM

MACRO AN4M12HM
    CLASS CORE ;
    FOREIGN AN4M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.398  LAYER ME1  ;
        ANTENNAGATEAREA 0.398  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.723  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.130 1.100 1.330 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.520 1.080 1.520 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.398  LAYER ME1  ;
        ANTENNAGATEAREA 0.398  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.723  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.080 1.080 3.080 1.400 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.980 1.540 9.260 2.100 ;
        RECT  6.940 0.680 9.220 0.880 ;
        RECT  9.020 0.410 9.220 0.880 ;
        RECT  6.900 1.540 9.260 1.740 ;
        RECT  7.790 0.680 8.390 1.740 ;
        RECT  7.940 0.680 8.220 2.100 ;
        RECT  7.980 0.410 8.180 2.100 ;
        RECT  6.900 1.540 7.180 2.100 ;
        RECT  6.940 0.410 7.140 0.880 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.398  LAYER ME1  ;
        ANTENNAGATEAREA 0.398  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.723  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.130 4.300 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.400 ;
        LAYER ME1 ;
        RECT  3.640 1.080 4.640 1.400 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.398  LAYER ME1  ;
        ANTENNAGATEAREA 0.398  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.723  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  5.700 1.130 5.900 1.330 ;
        LAYER ME2 ;
        RECT  5.700 0.840 5.900 1.400 ;
        LAYER ME1 ;
        RECT  5.200 1.080 6.200 1.400 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 10.000 2.540 ;
        RECT  9.500 1.540 9.780 2.540 ;
        RECT  8.460 1.900 8.740 2.540 ;
        RECT  7.420 1.900 7.700 2.540 ;
        RECT  6.360 1.900 6.640 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.710 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 10.000 0.140 ;
        RECT  9.540 -0.140 9.740 0.690 ;
        RECT  8.460 -0.140 8.740 0.520 ;
        RECT  7.420 -0.140 7.700 0.520 ;
        RECT  6.400 -0.140 6.600 0.710 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.300 2.980 0.460 ;
        RECT  0.620 0.300 0.900 0.520 ;
        RECT  1.660 0.300 1.940 0.520 ;
        RECT  2.700 0.300 2.980 0.520 ;
        RECT  3.220 0.300 3.500 0.880 ;
        RECT  2.170 0.680 4.540 0.880 ;
        RECT  3.740 0.300 5.000 0.460 ;
        RECT  3.740 0.300 4.020 0.520 ;
        RECT  4.780 0.300 5.000 0.880 ;
        RECT  5.860 0.430 6.060 0.880 ;
        RECT  4.780 0.680 6.060 0.880 ;
        RECT  0.140 0.430 0.340 0.880 ;
        RECT  0.140 0.680 1.900 0.880 ;
        RECT  6.540 1.080 7.590 1.280 ;
        RECT  6.540 1.080 6.740 1.740 ;
        RECT  0.660 1.580 6.740 1.740 ;
        RECT  0.660 1.580 0.860 1.990 ;
        RECT  1.700 0.680 1.900 1.990 ;
        RECT  2.740 1.580 2.940 1.990 ;
        RECT  3.780 1.580 3.980 1.990 ;
        RECT  4.820 1.580 5.020 1.990 ;
        RECT  5.860 1.580 6.060 1.990 ;
        RECT  8.570 1.080 9.320 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.470 2.400 ;
        RECT  6.250 1.140 10.000 2.400 ;
        RECT  0.000 1.290 10.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 10.000 1.140 ;
        RECT  0.470 0.000 6.250 1.290 ;
    END
END AN4M12HM

MACRO AN4M0HM
    CLASS CORE ;
    FOREIGN AN4M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        ANTENNAGATEAREA 0.080  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 5.045  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.130 1.900 1.330 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.560 ;
        LAYER ME1 ;
        RECT  1.700 1.040 2.100 1.420 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.400 0.840 0.700 1.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.100 1.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.080  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.300 0.840 1.540 1.400 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.700 1.880 3.100 2.080 ;
        RECT  2.900 0.330 3.100 2.080 ;
        RECT  2.700 0.330 3.100 0.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.840 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.100 -0.140 2.380 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 0.440 1.940 0.640 ;
        RECT  1.740 0.440 1.940 0.860 ;
        RECT  1.740 0.660 2.540 0.860 ;
        RECT  2.340 0.660 2.540 1.740 ;
        RECT  0.620 1.580 2.540 1.740 ;
        RECT  0.620 1.580 0.900 2.100 ;
        RECT  1.660 1.580 1.940 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AN4M0HM

MACRO AN3M8HM
    CLASS CORE ;
    FOREIGN AN3M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.241  LAYER ME1  ;
        ANTENNAGATEAREA 0.241  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.919  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.700 1.080 1.900 1.280 ;
        LAYER ME2 ;
        RECT  1.700 0.840 1.900 1.400 ;
        LAYER ME1 ;
        RECT  1.560 1.080 2.250 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.241  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 0.660 2.800 1.280 ;
        RECT  0.960 0.660 2.800 0.860 ;
        RECT  0.960 0.660 1.240 1.280 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.241  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.440 3.260 1.600 ;
        RECT  3.060 1.020 3.260 1.600 ;
        RECT  0.500 1.020 0.700 1.600 ;
        END
    END C
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.020 0.660 5.300 2.100 ;
        RECT  5.060 0.390 5.300 2.100 ;
        RECT  3.980 1.540 5.300 1.720 ;
        RECT  4.900 0.660 5.300 1.720 ;
        RECT  4.020 0.660 5.300 0.860 ;
        RECT  3.980 1.540 4.260 2.100 ;
        RECT  4.020 0.390 4.220 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.580 1.480 5.780 2.540 ;
        RECT  4.500 1.900 4.780 2.540 ;
        RECT  3.420 2.080 3.700 2.540 ;
        RECT  2.300 2.080 2.580 2.540 ;
        RECT  1.180 2.080 1.460 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.580 -0.140 5.780 0.660 ;
        RECT  4.500 -0.140 4.780 0.500 ;
        RECT  3.320 -0.140 3.600 0.540 ;
        RECT  0.340 -0.140 0.540 0.670 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.700 0.340 3.160 0.500 ;
        RECT  3.000 0.340 3.160 0.860 ;
        RECT  3.000 0.700 3.820 0.860 ;
        RECT  3.660 1.020 4.700 1.220 ;
        RECT  3.660 0.700 3.820 1.920 ;
        RECT  0.580 1.760 3.820 1.920 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END AN3M8HM

MACRO AN3M6HM
    CLASS CORE ;
    FOREIGN AN3M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.220 0.660 3.500 2.100 ;
        RECT  3.260 0.390 3.500 2.100 ;
        RECT  2.180 1.540 3.500 1.720 ;
        RECT  2.220 0.660 3.500 0.860 ;
        RECT  2.180 1.540 2.460 2.100 ;
        RECT  2.220 0.390 2.420 0.860 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        ANTENNAGATEAREA 0.134  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.863  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.140 1.500 1.340 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.080 1.700 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.420 1.300 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.134  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 0.840 1.100 1.330 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.600 0.140 ;
        RECT  2.700 -0.140 2.980 0.500 ;
        RECT  1.720 -0.140 1.920 0.580 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.600 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    OBS
        LAYER ME1 ;
        RECT  0.100 0.340 1.500 0.540 ;
        RECT  1.340 0.340 1.500 0.900 ;
        RECT  1.340 0.740 2.020 0.900 ;
        RECT  1.860 1.020 2.760 1.220 ;
        RECT  1.860 0.740 2.020 1.740 ;
        RECT  0.100 1.580 2.020 1.740 ;
        RECT  1.100 1.580 1.460 1.780 ;
        RECT  0.100 1.580 0.420 1.800 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.600 1.140 ;
    END
END AN3M6HM

MACRO AN3M4HM
    CLASS CORE ;
    FOREIGN AN3M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        ANTENNAGATEAREA 0.122  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.314  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.040 1.700 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.440 0.840 0.700 1.420 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.122  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 0.840 1.140 1.400 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.300 1.540 3.100 1.740 ;
        RECT  2.900 0.660 3.100 1.740 ;
        RECT  2.340 0.660 3.100 0.860 ;
        RECT  2.300 1.540 2.580 2.100 ;
        RECT  2.340 0.390 2.540 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.820 1.900 3.100 2.540 ;
        RECT  1.780 1.900 2.060 2.540 ;
        RECT  0.740 1.900 1.020 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.820 -0.140 3.100 0.500 ;
        RECT  1.700 -0.140 1.980 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 0.360 1.540 0.560 ;
        RECT  1.340 0.360 1.540 0.860 ;
        RECT  1.340 0.660 2.140 0.860 ;
        RECT  1.940 1.040 2.740 1.320 ;
        RECT  1.940 0.660 2.140 1.740 ;
        RECT  0.260 1.580 2.140 1.740 ;
        RECT  0.260 1.580 0.460 2.040 ;
        RECT  1.300 1.580 1.500 2.040 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AN3M4HM

MACRO AN3M2HM
    CLASS CORE ;
    FOREIGN AN3M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.040 1.600 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.830 0.540 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.830 1.100 1.400 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.240 1.440 2.700 2.080 ;
        RECT  2.500 0.330 2.700 2.080 ;
        RECT  2.200 0.330 2.700 0.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.680 1.900 1.960 2.540 ;
        RECT  0.640 1.900 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.620 -0.140 1.900 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.430 1.460 0.630 ;
        RECT  1.260 0.430 1.460 0.860 ;
        RECT  1.260 0.660 2.060 0.860 ;
        RECT  1.860 0.660 2.060 1.740 ;
        RECT  0.120 1.580 2.060 1.740 ;
        RECT  0.120 1.580 0.400 2.100 ;
        RECT  1.160 1.580 1.440 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AN3M2HM

MACRO AN3M1HM
    CLASS CORE ;
    FOREIGN AN3M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.040 1.600 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.830 0.540 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.840 1.100 1.370 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 1.880 2.700 2.080 ;
        RECT  2.500 0.350 2.700 2.080 ;
        RECT  2.200 0.350 2.700 0.550 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.680 1.900 1.960 2.540 ;
        RECT  0.640 1.900 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.600 -0.140 1.880 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.430 1.440 0.630 ;
        RECT  1.260 0.430 1.440 0.860 ;
        RECT  1.260 0.660 2.040 0.860 ;
        RECT  1.840 0.660 2.040 1.740 ;
        RECT  0.120 1.580 2.040 1.740 ;
        RECT  0.120 1.580 0.400 2.100 ;
        RECT  1.160 1.580 1.440 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AN3M1HM

MACRO AN3M16HM
    CLASS CORE ;
    FOREIGN AN3M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.130 1.100 1.330 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.500 1.080 1.540 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.060 1.080 3.100 1.360 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.420 1.540 8.700 2.060 ;
        RECT  5.340 0.680 8.660 0.880 ;
        RECT  8.460 0.410 8.660 0.880 ;
        RECT  5.300 1.540 8.700 1.740 ;
        RECT  7.380 1.540 7.660 2.060 ;
        RECT  7.420 0.410 7.620 0.880 ;
        RECT  6.900 0.680 7.500 1.740 ;
        RECT  6.340 1.540 6.620 2.060 ;
        RECT  6.380 0.410 6.580 0.880 ;
        RECT  5.300 1.540 5.580 2.060 ;
        RECT  5.340 0.410 5.540 0.880 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.426  LAYER ME1  ;
        ANTENNAGATEAREA 0.426  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.685  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.130 4.300 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.400 ;
        LAYER ME1 ;
        RECT  3.600 1.080 4.700 1.360 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.940 1.540 9.220 2.540 ;
        RECT  7.900 1.900 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.980 -0.140 9.180 0.690 ;
        RECT  7.900 -0.140 8.180 0.520 ;
        RECT  6.860 -0.140 7.140 0.520 ;
        RECT  5.820 -0.140 6.100 0.520 ;
        RECT  4.820 -0.140 5.020 0.710 ;
        RECT  3.740 -0.140 4.020 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.300 2.980 0.460 ;
        RECT  0.620 0.300 0.900 0.520 ;
        RECT  1.660 0.300 1.940 0.520 ;
        RECT  2.700 0.300 2.980 0.520 ;
        RECT  2.180 0.620 2.460 0.880 ;
        RECT  3.260 0.480 3.460 0.880 ;
        RECT  4.300 0.480 4.500 0.880 ;
        RECT  2.180 0.680 4.500 0.880 ;
        RECT  0.140 0.430 0.340 0.880 ;
        RECT  1.140 0.620 1.420 0.880 ;
        RECT  0.140 0.680 1.900 0.880 ;
        RECT  4.900 1.080 6.700 1.280 ;
        RECT  1.700 0.680 1.900 1.740 ;
        RECT  4.900 1.080 5.100 1.740 ;
        RECT  0.140 1.540 5.100 1.740 ;
        RECT  0.140 1.540 0.340 2.030 ;
        RECT  1.180 1.540 1.380 2.030 ;
        RECT  2.220 1.540 2.420 2.030 ;
        RECT  3.260 1.540 3.460 2.030 ;
        RECT  4.300 1.540 4.500 2.030 ;
        RECT  7.700 1.080 8.780 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.460 2.400 ;
        RECT  4.660 1.140 9.600 2.400 ;
        RECT  0.000 1.290 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
        RECT  0.460 0.000 4.660 1.290 ;
    END
END AN3M16HM

MACRO AN3M12HM
    CLASS CORE ;
    FOREIGN AN3M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.373  LAYER ME1  ;
        ANTENNAGATEAREA 0.373  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.839  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.130 1.100 1.330 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.500 1.080 1.540 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.373  LAYER ME1  ;
        ANTENNAGATEAREA 0.373  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.839  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.060 1.080 3.100 1.360 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  7.380 1.540 7.660 2.060 ;
        RECT  5.340 0.680 7.620 0.880 ;
        RECT  7.420 0.410 7.620 0.880 ;
        RECT  5.300 1.540 7.660 1.740 ;
        RECT  6.100 0.680 6.700 1.740 ;
        RECT  6.340 0.680 6.620 2.060 ;
        RECT  6.380 0.410 6.580 2.060 ;
        RECT  5.300 1.540 5.580 2.060 ;
        RECT  5.340 0.410 5.540 0.880 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.373  LAYER ME1  ;
        ANTENNAGATEAREA 0.373  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.923  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.100 1.130 4.300 1.330 ;
        LAYER ME2 ;
        RECT  4.100 0.840 4.300 1.400 ;
        LAYER ME1 ;
        RECT  3.600 1.080 4.700 1.360 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.400 2.540 ;
        RECT  7.900 1.540 8.180 2.540 ;
        RECT  6.860 1.900 7.140 2.540 ;
        RECT  5.820 1.900 6.100 2.540 ;
        RECT  4.780 1.900 5.060 2.540 ;
        RECT  3.740 1.900 4.020 2.540 ;
        RECT  2.700 1.900 2.980 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.400 0.140 ;
        RECT  7.940 -0.140 8.140 0.710 ;
        RECT  6.860 -0.140 7.140 0.520 ;
        RECT  5.820 -0.140 6.100 0.520 ;
        RECT  4.820 -0.140 5.020 0.710 ;
        RECT  3.740 -0.140 4.020 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.300 2.980 0.460 ;
        RECT  0.620 0.300 0.900 0.520 ;
        RECT  1.660 0.300 1.940 0.520 ;
        RECT  2.700 0.300 2.980 0.520 ;
        RECT  2.180 0.620 2.460 0.880 ;
        RECT  3.260 0.480 3.460 0.880 ;
        RECT  4.300 0.480 4.500 0.880 ;
        RECT  2.180 0.680 4.500 0.880 ;
        RECT  0.140 0.430 0.340 0.880 ;
        RECT  1.140 0.620 1.420 0.880 ;
        RECT  0.140 0.680 1.900 0.880 ;
        RECT  4.900 1.080 5.900 1.280 ;
        RECT  1.700 0.680 1.900 1.740 ;
        RECT  4.900 1.080 5.100 1.740 ;
        RECT  0.140 1.540 5.100 1.740 ;
        RECT  0.140 1.540 0.340 2.030 ;
        RECT  1.180 1.540 1.380 2.030 ;
        RECT  2.220 1.540 2.420 2.030 ;
        RECT  3.260 1.540 3.460 2.030 ;
        RECT  4.300 1.540 4.500 2.030 ;
        RECT  6.990 1.080 7.710 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.460 2.400 ;
        RECT  4.660 1.140 8.400 2.400 ;
        RECT  0.000 1.290 8.400 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.400 1.140 ;
        RECT  0.460 0.000 4.660 1.290 ;
    END
END AN3M12HM

MACRO AN3M0HM
    CLASS CORE ;
    FOREIGN AN3M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        ANTENNAGATEAREA 0.076  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 4.677  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.130 1.500 1.330 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.560 ;
        LAYER ME1 ;
        RECT  1.300 1.040 1.600 1.420 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.830 0.600 1.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.076  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.800 0.830 1.100 1.400 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.200 1.880 2.700 2.080 ;
        RECT  2.500 0.310 2.700 2.080 ;
        RECT  2.260 0.310 2.700 0.660 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  1.680 1.900 1.960 2.540 ;
        RECT  0.640 1.900 0.920 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  1.600 -0.140 1.880 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.100 0.430 1.440 0.630 ;
        RECT  1.260 0.430 1.440 0.860 ;
        RECT  1.260 0.660 2.060 0.860 ;
        RECT  1.860 0.660 2.060 1.740 ;
        RECT  0.120 1.580 2.060 1.740 ;
        RECT  0.120 1.580 0.400 2.100 ;
        RECT  1.160 1.580 1.440 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AN3M0HM

MACRO AN2M8HM
    CLASS CORE ;
    FOREIGN AN2M8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        ANTENNAGATEAREA 0.230  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.167  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  1.300 1.080 1.500 1.280 ;
        LAYER ME2 ;
        RECT  1.300 0.840 1.500 1.400 ;
        LAYER ME1 ;
        RECT  0.900 1.020 1.540 1.340 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.230  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.120 2.120 1.340 ;
        RECT  1.700 0.660 1.900 1.340 ;
        RECT  0.500 0.660 1.900 0.860 ;
        RECT  0.500 0.660 0.700 1.340 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.880 1.540 4.160 2.100 ;
        RECT  2.880 0.660 4.160 0.860 ;
        RECT  3.920 0.390 4.160 0.860 ;
        RECT  3.700 0.660 3.920 1.740 ;
        RECT  2.840 1.540 4.160 1.740 ;
        RECT  2.840 1.540 3.120 2.100 ;
        RECT  2.880 0.390 3.080 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.800 2.540 ;
        RECT  4.400 1.450 4.680 2.540 ;
        RECT  3.360 1.900 3.640 2.540 ;
        RECT  2.250 1.860 2.530 2.540 ;
        RECT  1.140 1.860 1.420 2.540 ;
        RECT  0.140 1.750 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.800 0.140 ;
        RECT  4.400 -0.140 4.680 0.720 ;
        RECT  3.360 -0.140 3.640 0.500 ;
        RECT  2.380 -0.140 2.580 0.600 ;
        RECT  0.300 -0.140 0.580 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  1.100 0.340 2.220 0.500 ;
        RECT  2.060 0.340 2.220 0.940 ;
        RECT  2.060 0.760 2.680 0.940 ;
        RECT  2.520 1.020 3.500 1.220 ;
        RECT  2.520 0.760 2.680 1.700 ;
        RECT  0.660 1.540 2.680 1.700 ;
        RECT  0.660 1.540 0.860 2.030 ;
        RECT  1.700 1.540 1.900 2.030 ;
        LAYER VTPH ;
        RECT  0.000 1.140 4.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 4.800 1.140 ;
    END
END AN2M8HM

MACRO AN2M6HM
    CLASS CORE ;
    FOREIGN AN2M6HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        ANTENNAGATEAREA 0.149  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 3.565  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.160 1.100 1.360 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.560 ;
        LAYER ME1 ;
        RECT  0.500 1.060 1.200 1.380 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.149  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.980 0.320 1.600 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.740 1.540 3.100 2.100 ;
        RECT  2.900 0.390 3.100 2.100 ;
        RECT  1.740 0.660 3.100 0.860 ;
        RECT  2.780 0.390 3.100 0.860 ;
        RECT  1.700 1.540 3.100 1.720 ;
        RECT  1.700 1.540 1.980 2.100 ;
        RECT  1.740 0.390 1.940 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 3.200 2.540 ;
        RECT  2.220 1.900 2.500 2.540 ;
        RECT  1.180 1.860 1.460 2.540 ;
        RECT  0.100 1.880 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 3.200 0.140 ;
        RECT  2.220 -0.140 2.500 0.500 ;
        RECT  1.160 -0.140 1.360 0.580 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.380 1.000 0.580 ;
        RECT  0.840 0.380 1.000 0.900 ;
        RECT  0.840 0.740 1.520 0.900 ;
        RECT  1.360 1.020 2.520 1.220 ;
        RECT  1.360 0.740 1.520 1.700 ;
        RECT  0.660 1.540 1.520 1.700 ;
        RECT  0.660 1.540 0.940 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 3.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 3.200 1.140 ;
    END
END AN2M6HM

MACRO AN2M4HM
    CLASS CORE ;
    FOREIGN AN2M4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.500 1.080 0.740 1.690 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.119  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.900 1.080 1.400 1.280 ;
        RECT  0.900 0.840 1.100 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.940 1.540 2.700 1.740 ;
        RECT  2.500 0.660 2.700 1.740 ;
        RECT  1.940 0.660 2.700 0.860 ;
        RECT  1.940 1.540 2.140 1.920 ;
        RECT  1.940 0.430 2.140 0.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.800 2.540 ;
        RECT  2.420 1.900 2.700 2.540 ;
        RECT  1.380 1.860 1.660 2.540 ;
        RECT  0.300 1.850 0.580 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.800 0.140 ;
        RECT  2.420 -0.140 2.700 0.500 ;
        RECT  1.340 -0.140 1.620 0.360 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.420 0.520 1.720 0.680 ;
        RECT  1.560 1.040 2.300 1.320 ;
        RECT  1.560 0.520 1.720 1.700 ;
        RECT  0.900 1.540 1.720 1.700 ;
        RECT  0.900 1.540 1.100 2.020 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.800 1.140 ;
    END
END AN2M4HM

MACRO AN2M2HM
    CLASS CORE ;
    FOREIGN AN2M2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.520 1.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.280 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.390 1.900 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.100 2.020 1.300 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.040 -0.140 1.320 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.140 0.310 0.340 0.660 ;
        RECT  0.140 0.480 1.520 0.660 ;
        RECT  1.320 0.480 1.520 1.680 ;
        RECT  0.620 1.480 1.520 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END AN2M2HM

MACRO AN2M1HM
    CLASS CORE ;
    FOREIGN AN2M1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.600 1.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.220 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.390 1.900 1.790 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.100 2.020 1.300 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.040 -0.140 1.320 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 0.380 0.380 0.660 ;
        RECT  0.180 0.480 1.520 0.660 ;
        RECT  1.320 0.480 1.520 1.680 ;
        RECT  0.620 1.480 1.520 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END AN2M1HM

MACRO AN2M16HM
    CLASS CORE ;
    FOREIGN AN2M16HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.406  LAYER ME1  ;
        ANTENNAGATEAREA 0.406  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.692  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.130 1.100 1.330 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.500 1.080 1.540 1.360 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.406  LAYER ME1  ;
        ANTENNAGATEAREA 0.406  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.769  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.040 1.080 3.140 1.360 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.984  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.860 1.540 7.140 2.060 ;
        RECT  3.780 0.680 7.100 0.880 ;
        RECT  6.900 0.410 7.100 0.880 ;
        RECT  3.740 1.540 7.140 1.740 ;
        RECT  5.820 1.540 6.100 2.060 ;
        RECT  5.860 0.410 6.060 0.880 ;
        RECT  5.300 0.680 5.600 1.740 ;
        RECT  4.780 1.540 5.060 2.060 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  3.740 1.540 4.020 2.060 ;
        RECT  3.780 0.410 3.980 0.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 8.000 2.540 ;
        RECT  7.380 1.540 7.660 2.540 ;
        RECT  6.340 1.900 6.620 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 8.000 0.140 ;
        RECT  7.380 -0.140 7.660 0.520 ;
        RECT  6.340 -0.140 6.620 0.520 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.260 -0.140 3.460 0.710 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.620 0.900 0.880 ;
        RECT  1.700 0.480 1.900 0.880 ;
        RECT  2.740 0.480 2.940 0.880 ;
        RECT  0.620 0.680 2.940 0.880 ;
        RECT  0.140 0.300 1.420 0.460 ;
        RECT  1.140 0.300 1.420 0.520 ;
        RECT  3.340 1.080 5.140 1.280 ;
        RECT  0.140 0.300 0.340 1.740 ;
        RECT  3.340 1.080 3.540 1.740 ;
        RECT  0.140 1.540 3.540 1.740 ;
        RECT  0.660 1.540 0.860 2.030 ;
        RECT  1.700 1.540 1.900 2.030 ;
        RECT  2.740 1.540 2.940 2.030 ;
        RECT  5.880 1.080 7.320 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.460 2.400 ;
        RECT  3.100 1.140 8.000 2.400 ;
        RECT  0.000 1.250 8.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 8.000 1.140 ;
        RECT  0.460 0.000 3.100 1.250 ;
    END
END AN2M16HM

MACRO AN2M12HM
    CLASS CORE ;
    FOREIGN AN2M12HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.352  LAYER ME1  ;
        ANTENNAGATEAREA 0.352  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 1.952  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.900 1.130 1.100 1.330 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.100 1.400 ;
        LAYER ME1 ;
        RECT  0.500 1.080 1.540 1.360 ;
        END
    END A
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.488  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.820 1.540 6.100 2.060 ;
        RECT  3.780 0.680 6.060 0.880 ;
        RECT  5.860 0.410 6.060 0.880 ;
        RECT  3.740 1.540 6.100 1.740 ;
        RECT  4.780 1.540 5.060 2.060 ;
        RECT  4.820 0.410 5.020 0.880 ;
        RECT  4.500 0.680 4.760 1.740 ;
        RECT  3.740 1.540 4.020 2.060 ;
        RECT  3.780 0.410 3.980 0.880 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.352  LAYER ME1  ;
        ANTENNAGATEAREA 0.352  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 2.041  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  2.500 1.130 2.700 1.330 ;
        LAYER ME2 ;
        RECT  2.500 0.840 2.700 1.400 ;
        LAYER ME1 ;
        RECT  2.040 1.080 3.140 1.360 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.800 2.540 ;
        RECT  6.380 1.480 6.580 2.540 ;
        RECT  5.300 1.900 5.580 2.540 ;
        RECT  4.260 1.900 4.540 2.540 ;
        RECT  3.220 1.900 3.500 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.800 0.140 ;
        RECT  6.380 -0.140 6.580 0.690 ;
        RECT  5.300 -0.140 5.580 0.520 ;
        RECT  4.260 -0.140 4.540 0.520 ;
        RECT  3.260 -0.140 3.460 0.710 ;
        RECT  2.180 -0.140 2.460 0.520 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.620 0.620 0.900 0.880 ;
        RECT  1.700 0.410 1.900 0.880 ;
        RECT  2.740 0.480 2.940 0.880 ;
        RECT  0.620 0.680 2.940 0.880 ;
        RECT  0.140 0.300 1.420 0.460 ;
        RECT  1.140 0.300 1.420 0.520 ;
        RECT  3.340 1.080 4.340 1.280 ;
        RECT  0.140 0.300 0.340 1.740 ;
        RECT  3.340 1.080 3.540 1.740 ;
        RECT  0.140 1.540 3.540 1.740 ;
        RECT  0.660 1.540 0.860 2.030 ;
        RECT  1.700 1.540 1.900 2.030 ;
        RECT  2.740 1.540 2.940 2.030 ;
        RECT  5.340 1.080 6.050 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 0.460 2.400 ;
        RECT  3.100 1.140 6.800 2.400 ;
        RECT  0.000 1.250 6.800 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 6.800 1.140 ;
        RECT  0.460 0.000 3.100 1.250 ;
    END
END AN2M12HM

MACRO AN2M0HM
    CLASS CORE ;
    FOREIGN AN2M0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.840 0.600 1.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.071  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.860 0.840 1.140 1.240 ;
        END
    END B
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.680 0.390 1.900 1.770 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 2.000 2.540 ;
        RECT  1.100 2.020 1.300 2.540 ;
        RECT  0.100 1.500 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 2.000 0.140 ;
        RECT  1.040 -0.140 1.320 0.320 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.180 0.380 0.380 0.660 ;
        RECT  0.180 0.480 1.520 0.660 ;
        RECT  1.320 0.480 1.520 1.680 ;
        RECT  0.620 1.480 1.520 1.680 ;
        LAYER VTPH ;
        RECT  0.000 1.140 2.000 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 2.000 1.140 ;
    END
END AN2M0HM

MACRO ADHM8HM
    CLASS CORE ;
    FOREIGN ADHM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.312  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.260 1.120 5.700 1.560 ;
        RECT  3.170 1.120 5.700 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.312  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.440 1.440 4.560 1.600 ;
        RECT  2.440 1.180 3.000 1.600 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.700 1.470 1.900 1.980 ;
        RECT  0.660 0.680 1.900 0.840 ;
        RECT  1.700 0.370 1.900 0.840 ;
        RECT  0.660 1.470 1.900 1.670 ;
        RECT  1.300 0.680 1.500 1.670 ;
        RECT  0.660 1.470 0.860 1.980 ;
        RECT  0.660 0.370 0.860 0.840 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.944  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  8.420 1.470 8.620 1.970 ;
        RECT  7.380 0.660 8.620 0.840 ;
        RECT  8.420 0.370 8.620 0.840 ;
        RECT  7.380 1.470 8.620 1.670 ;
        RECT  7.700 0.660 7.900 1.670 ;
        RECT  7.380 1.470 7.580 1.970 ;
        RECT  7.380 0.370 7.580 0.840 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 9.600 2.540 ;
        RECT  8.900 1.900 9.180 2.540 ;
        RECT  7.860 1.900 8.140 2.540 ;
        RECT  6.860 1.470 7.060 2.540 ;
        RECT  6.380 1.840 6.580 2.540 ;
        RECT  4.460 1.810 4.660 2.540 ;
        RECT  3.340 2.080 3.620 2.540 ;
        RECT  2.220 2.080 2.500 2.540 ;
        RECT  1.140 1.900 1.420 2.540 ;
        RECT  0.140 1.480 0.340 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 9.600 0.140 ;
        RECT  8.900 -0.140 9.180 0.500 ;
        RECT  7.860 -0.140 8.140 0.500 ;
        RECT  6.860 -0.140 7.060 0.650 ;
        RECT  5.260 -0.140 5.540 0.320 ;
        RECT  4.260 -0.140 4.460 0.580 ;
        RECT  2.360 -0.140 2.560 0.580 ;
        RECT  1.140 -0.140 1.420 0.500 ;
        RECT  0.140 -0.140 0.340 0.650 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.460 1.000 1.100 1.280 ;
        RECT  4.660 0.480 6.140 0.640 ;
        RECT  3.380 0.300 3.580 0.960 ;
        RECT  2.090 0.800 6.220 0.960 ;
        RECT  1.700 1.040 2.250 1.240 ;
        RECT  6.020 0.800 6.220 1.280 ;
        RECT  2.090 0.800 2.250 1.920 ;
        RECT  2.090 1.760 4.140 1.920 ;
        RECT  2.820 1.760 3.020 2.100 ;
        RECT  3.940 1.760 4.140 2.100 ;
        RECT  6.380 1.040 7.500 1.240 ;
        RECT  6.380 0.360 6.580 1.630 ;
        RECT  5.860 1.470 6.580 1.630 ;
        RECT  5.860 1.470 6.060 2.060 ;
        RECT  8.100 1.000 8.740 1.280 ;
        LAYER VTPH ;
        RECT  0.000 1.140 9.600 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 9.600 1.140 ;
    END
END ADHM8HM

MACRO ADHM4HM
    CLASS CORE ;
    FOREIGN ADHM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.100 1.120 4.660 1.560 ;
        RECT  2.130 1.120 4.660 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.540 1.440 3.520 1.600 ;
        RECT  1.540 1.180 1.960 1.600 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.660 1.470 0.860 1.980 ;
        RECT  0.100 0.680 0.860 0.840 ;
        RECT  0.660 0.370 0.860 0.840 ;
        RECT  0.100 1.470 0.860 1.670 ;
        RECT  0.100 0.680 0.300 1.670 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  6.340 1.470 7.100 1.670 ;
        RECT  6.900 0.660 7.100 1.670 ;
        RECT  6.340 0.660 7.100 0.840 ;
        RECT  6.340 1.470 6.540 1.970 ;
        RECT  6.340 0.370 6.540 0.840 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 7.200 2.540 ;
        RECT  6.820 1.900 7.100 2.540 ;
        RECT  5.820 1.470 6.020 2.540 ;
        RECT  5.340 1.840 5.540 2.540 ;
        RECT  3.420 1.810 3.620 2.540 ;
        RECT  2.300 2.080 2.580 2.540 ;
        RECT  1.180 2.080 1.460 2.540 ;
        RECT  0.100 1.900 0.380 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 7.200 0.140 ;
        RECT  6.820 -0.140 7.100 0.500 ;
        RECT  5.820 -0.140 6.020 0.650 ;
        RECT  4.220 -0.140 4.500 0.320 ;
        RECT  3.220 -0.140 3.420 0.580 ;
        RECT  1.320 -0.140 1.520 0.580 ;
        RECT  0.100 -0.140 0.380 0.500 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  3.620 0.480 5.100 0.640 ;
        RECT  2.340 0.300 2.540 0.960 ;
        RECT  1.050 0.800 5.180 0.960 ;
        RECT  0.660 1.040 1.210 1.240 ;
        RECT  4.980 0.800 5.180 1.280 ;
        RECT  1.050 0.800 1.210 1.920 ;
        RECT  1.050 1.760 3.100 1.920 ;
        RECT  1.780 1.760 1.980 2.100 ;
        RECT  2.900 1.760 3.100 2.100 ;
        RECT  5.340 1.040 6.580 1.240 ;
        RECT  5.340 0.360 5.540 1.630 ;
        RECT  4.820 1.470 5.540 1.630 ;
        RECT  4.820 1.470 5.020 2.060 ;
        LAYER VTPH ;
        RECT  0.000 1.140 7.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 7.200 1.140 ;
    END
END ADHM4HM

MACRO ADHM2HM
    CLASS CORE ;
    FOREIGN ADHM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER ME1  ;
        ANTENNAGATEAREA 0.175  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.203  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.160 1.140 1.360 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.140 2.680 1.300 ;
        RECT  0.840 1.140 1.230 1.390 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 1.460 3.120 1.670 ;
        RECT  2.840 1.140 3.120 1.670 ;
        END
    END A
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.410 0.320 2.100 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.700 1.440 5.100 2.100 ;
        RECT  4.900 0.450 5.100 2.100 ;
        RECT  4.700 0.450 5.100 0.650 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.220 1.440 4.420 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.220 -0.140 4.420 0.690 ;
        RECT  2.620 -0.140 2.900 0.340 ;
        RECT  0.720 -0.140 0.920 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.100 0.300 2.300 0.660 ;
        RECT  3.220 0.300 3.420 0.660 ;
        RECT  2.100 0.500 3.420 0.660 ;
        RECT  1.620 0.340 1.820 0.980 ;
        RECT  0.500 0.820 3.580 0.980 ;
        RECT  3.380 0.820 3.580 1.320 ;
        RECT  0.500 0.820 0.660 1.740 ;
        RECT  0.500 1.580 1.220 1.740 ;
        RECT  1.060 1.580 1.220 2.100 ;
        RECT  1.060 1.900 1.430 2.100 ;
        RECT  3.740 1.080 4.640 1.280 ;
        RECT  3.740 0.300 3.940 2.080 ;
        RECT  3.020 1.880 3.940 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END ADHM2HM

MACRO ADHM1HM
    CLASS CORE ;
    FOREIGN ADHM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME2  ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        ANTENNAMAXSIDEAREACAR 6.611  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.160 1.140 1.360 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.140 2.680 1.300 ;
        RECT  0.840 1.140 1.230 1.390 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.164  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 1.460 3.120 1.670 ;
        RECT  2.840 1.140 3.120 1.670 ;
        END
    END A
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.390 0.320 2.100 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.700 1.870 5.100 2.070 ;
        RECT  4.900 0.450 5.100 2.070 ;
        RECT  4.700 0.450 5.100 0.650 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.220 1.820 4.420 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.220 -0.140 4.420 0.690 ;
        RECT  2.620 -0.140 2.900 0.340 ;
        RECT  0.720 -0.140 0.920 0.660 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.100 0.300 2.300 0.660 ;
        RECT  3.220 0.300 3.420 0.660 ;
        RECT  2.100 0.500 3.420 0.660 ;
        RECT  1.620 0.340 1.820 0.980 ;
        RECT  0.500 0.820 3.580 0.980 ;
        RECT  3.380 0.820 3.580 1.320 ;
        RECT  0.500 0.820 0.660 1.740 ;
        RECT  0.500 1.580 1.220 1.740 ;
        RECT  1.060 1.580 1.220 2.100 ;
        RECT  1.060 1.900 1.430 2.100 ;
        RECT  3.740 1.080 4.640 1.280 ;
        RECT  3.740 0.300 3.940 2.080 ;
        RECT  3.020 1.880 3.940 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END ADHM1HM

MACRO ADHM0HM
    CLASS CORE ;
    FOREIGN ADHM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY X Y ;
    SITE CORE_6T ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        ANTENNAGATEAREA 0.157  LAYER ME2  ;
        ANTENNAMAXSIDEAREACAR 6.913  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  0.940 1.160 1.140 1.360 ;
        LAYER ME2 ;
        RECT  0.900 0.840 1.160 1.560 ;
        LAYER ME1 ;
        RECT  0.840 1.140 2.680 1.300 ;
        RECT  0.840 1.140 1.230 1.390 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  1.400 1.460 3.120 1.670 ;
        RECT  2.840 1.140 3.120 1.670 ;
        END
    END A
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 0.310 0.320 2.100 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.700 1.870 5.100 2.070 ;
        RECT  4.900 0.390 5.100 2.070 ;
        RECT  4.700 0.390 5.100 0.590 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.220 1.750 4.420 2.540 ;
        RECT  2.180 1.900 2.460 2.540 ;
        RECT  1.660 1.900 1.940 2.540 ;
        RECT  0.620 1.900 0.900 2.540 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.220 -0.140 4.420 0.630 ;
        RECT  2.620 -0.140 2.900 0.340 ;
        RECT  0.720 -0.140 0.920 0.560 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  2.100 0.300 2.300 0.660 ;
        RECT  3.220 0.300 3.420 0.660 ;
        RECT  2.100 0.500 3.420 0.660 ;
        RECT  1.620 0.310 1.820 0.980 ;
        RECT  0.500 0.820 3.580 0.980 ;
        RECT  3.380 0.820 3.580 1.320 ;
        RECT  0.500 0.820 0.660 1.740 ;
        RECT  0.500 1.580 1.220 1.740 ;
        RECT  1.060 1.580 1.220 2.100 ;
        RECT  1.060 1.900 1.430 2.100 ;
        RECT  3.740 1.080 4.640 1.280 ;
        RECT  3.740 0.300 3.940 2.080 ;
        RECT  3.020 1.880 3.940 2.080 ;
        LAYER VTPH ;
        RECT  0.000 1.140 5.200 2.400 ;
        LAYER VTNH ;
        RECT  0.000 0.000 5.200 1.140 ;
    END
END ADHM0HM

MACRO ADFM8HM
    CLASS CORE ;
    FOREIGN ADFM8HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.517  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.760 1.120 3.400 1.280 ;
        RECT  2.900 1.120 3.100 1.560 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.520  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.900 3.540 3.640 3.740 ;
        RECT  2.100 3.940 3.100 4.140 ;
        RECT  2.900 3.540 3.100 4.140 ;
        RECT  2.100 3.700 2.300 4.140 ;
        RECT  1.340 3.700 2.300 3.900 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.382  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.540 3.300 2.740 3.780 ;
        RECT  0.480 3.300 2.740 3.500 ;
        RECT  0.480 3.300 0.680 3.860 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.140 0.420 5.340 2.100 ;
        RECT  4.100 1.320 5.340 1.520 ;
        RECT  4.900 0.660 5.340 1.520 ;
        RECT  4.100 0.660 5.340 0.820 ;
        RECT  4.100 1.320 4.300 2.100 ;
        RECT  4.100 0.420 4.300 0.820 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  5.140 2.700 5.340 4.380 ;
        RECT  4.120 3.940 5.340 4.140 ;
        RECT  4.900 3.200 5.340 4.140 ;
        RECT  4.120 3.200 5.340 3.400 ;
        RECT  4.120 3.940 4.320 4.380 ;
        RECT  4.120 2.700 4.320 3.400 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 6.000 2.540 ;
        RECT  5.660 1.460 5.860 3.340 ;
        RECT  4.620 1.740 4.820 3.040 ;
        RECT  3.600 1.760 3.800 3.060 ;
        RECT  3.260 2.140 3.800 2.540 ;
        RECT  1.500 2.140 1.780 2.540 ;
        RECT  1.180 2.260 1.460 2.820 ;
        RECT  0.100 2.260 0.380 3.080 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 6.000 0.140 ;
        RECT  5.660 -0.140 5.860 0.600 ;
        RECT  4.580 -0.140 4.860 0.500 ;
        RECT  3.540 -0.140 3.820 0.640 ;
        RECT  1.500 -0.140 1.780 0.320 ;
        RECT  0.000 4.660 6.000 4.940 ;
        RECT  5.660 4.200 5.860 4.940 ;
        RECT  4.580 4.300 4.860 4.940 ;
        RECT  3.600 4.240 3.800 4.940 ;
        RECT  1.180 4.380 1.460 4.940 ;
        RECT  0.140 4.190 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 4.060 1.800 4.220 ;
        RECT  1.640 4.060 1.800 4.460 ;
        RECT  1.640 4.300 2.120 4.460 ;
        RECT  0.660 4.060 0.860 4.470 ;
        RECT  0.580 2.980 2.180 3.140 ;
        RECT  0.100 1.500 2.740 1.660 ;
        RECT  0.100 1.500 0.380 2.040 ;
        RECT  0.140 0.300 1.310 0.460 ;
        RECT  1.150 0.300 1.310 0.640 ;
        RECT  1.150 0.480 3.340 0.640 ;
        RECT  0.140 0.300 0.340 0.680 ;
        RECT  2.340 2.920 3.440 3.080 ;
        RECT  3.280 2.920 3.440 3.380 ;
        RECT  3.280 3.220 3.960 3.380 ;
        RECT  3.800 3.590 4.740 3.750 ;
        RECT  3.800 3.220 3.960 4.080 ;
        RECT  3.280 3.920 3.960 4.080 ;
        RECT  3.280 3.920 3.440 4.460 ;
        RECT  2.340 4.300 3.440 4.460 ;
        RECT  0.620 0.620 0.900 0.960 ;
        RECT  0.620 0.800 3.860 0.960 ;
        RECT  3.700 1.000 4.740 1.160 ;
        RECT  3.700 0.800 3.860 1.600 ;
        RECT  3.260 1.440 3.860 1.600 ;
        RECT  3.260 1.440 3.420 1.980 ;
        RECT  0.580 1.820 3.420 1.980 ;
        RECT  2.300 1.820 2.580 2.100 ;
        LAYER VTPH ;
        RECT  0.000 1.140 6.000 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 6.000 4.800 ;
        RECT  0.000 0.000 6.000 1.140 ;
    END
END ADFM8HM

MACRO ADFM4HM
    CLASS CORE ;
    FOREIGN ADFM4HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.530  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 3.520 1.280 ;
        RECT  0.100 0.840 0.360 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.521  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.920 3.500 3.640 3.700 ;
        RECT  2.100 3.940 3.080 4.140 ;
        RECT  2.920 3.500 3.080 4.140 ;
        RECT  2.100 3.440 2.300 4.140 ;
        RECT  1.340 3.440 2.300 3.640 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.404  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.500 3.080 2.740 3.740 ;
        RECT  0.480 3.080 2.740 3.280 ;
        RECT  0.480 3.080 0.680 3.680 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.120 1.440 4.700 1.670 ;
        RECT  4.500 0.660 4.700 1.670 ;
        RECT  4.120 0.660 4.700 0.820 ;
        RECT  4.120 1.440 4.320 2.080 ;
        RECT  4.120 0.390 4.320 0.820 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  4.120 3.980 4.700 4.140 ;
        RECT  4.500 3.090 4.700 4.140 ;
        RECT  4.120 3.090 4.700 3.370 ;
        RECT  4.120 3.980 4.320 4.300 ;
        RECT  4.120 2.720 4.320 3.370 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 5.200 2.540 ;
        RECT  4.580 1.900 4.860 2.920 ;
        RECT  3.540 1.780 3.820 2.920 ;
        RECT  0.140 2.260 0.340 2.980 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 5.200 0.140 ;
        RECT  4.580 -0.140 4.860 0.500 ;
        RECT  3.580 -0.140 3.780 0.590 ;
        RECT  1.750 -0.140 2.030 0.320 ;
        RECT  0.000 4.660 5.200 4.940 ;
        RECT  4.580 4.300 4.860 4.940 ;
        RECT  3.580 4.240 3.780 4.940 ;
        RECT  1.220 4.220 1.420 4.940 ;
        RECT  0.140 4.130 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 3.840 1.940 4.000 ;
        RECT  0.660 3.840 0.860 4.460 ;
        RECT  1.740 3.840 1.940 4.460 ;
        RECT  0.580 2.760 2.180 2.920 ;
        RECT  0.140 1.450 2.800 1.610 ;
        RECT  0.140 1.450 0.340 1.860 ;
        RECT  0.140 0.300 1.530 0.460 ;
        RECT  1.370 0.300 1.530 0.640 ;
        RECT  1.370 0.480 3.340 0.640 ;
        RECT  0.140 0.300 0.340 0.650 ;
        RECT  0.660 0.620 0.940 0.960 ;
        RECT  0.660 0.800 3.960 0.960 ;
        RECT  3.800 0.990 4.170 1.190 ;
        RECT  3.800 0.800 3.960 1.620 ;
        RECT  3.190 1.460 3.960 1.620 ;
        RECT  3.190 1.460 3.350 1.990 ;
        RECT  0.580 1.770 3.350 1.990 ;
        RECT  2.340 2.760 3.260 2.920 ;
        RECT  3.100 2.760 3.260 3.240 ;
        RECT  3.100 3.080 3.960 3.240 ;
        RECT  3.800 3.570 4.180 3.770 ;
        RECT  3.800 3.080 3.960 4.020 ;
        RECT  3.240 3.860 3.960 4.020 ;
        RECT  3.240 3.860 3.400 4.460 ;
        RECT  2.340 4.300 3.400 4.460 ;
        LAYER VTPH ;
        RECT  2.270 1.090 3.000 3.660 ;
        RECT  0.000 1.140 5.200 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 5.200 4.800 ;
        RECT  0.000 0.000 5.200 1.090 ;
        RECT  0.000 0.000 2.270 1.140 ;
        RECT  3.000 0.000 5.200 1.140 ;
    END
END ADFM4HM

MACRO ADFM2HM
    CLASS CORE ;
    FOREIGN ADFM2HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER ME1  ;
        ANTENNADIFFAREA 0.422  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.010 4.200 4.210 4.400 ;
        LAYER ME2 ;
        RECT  3.910 4.000 4.300 4.400 ;
        LAYER ME1 ;
        RECT  3.910 4.200 4.300 4.500 ;
        RECT  4.130 2.750 4.300 4.500 ;
        RECT  3.970 2.750 4.300 2.960 ;
        END
    END S
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.422  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 3.400 1.280 ;
        RECT  0.100 0.840 0.360 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.414  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.830 3.520 3.590 3.680 ;
        RECT  2.010 3.980 2.990 4.140 ;
        RECT  2.830 3.520 2.990 4.140 ;
        RECT  2.010 3.460 2.300 4.140 ;
        RECT  1.340 3.460 2.300 3.640 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.306  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.490 3.130 2.650 3.780 ;
        RECT  0.480 3.130 2.650 3.290 ;
        RECT  0.480 3.130 0.700 3.680 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.418  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.980 0.390 4.300 2.080 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.450 2.260 3.730 2.970 ;
        RECT  3.420 1.780 3.700 2.540 ;
        RECT  0.140 2.260 0.340 2.980 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.460 -0.140 3.660 0.590 ;
        RECT  1.750 -0.140 2.030 0.320 ;
        RECT  0.000 4.660 4.400 4.940 ;
        RECT  3.490 4.240 3.690 4.940 ;
        RECT  1.180 4.220 1.380 4.940 ;
        RECT  0.140 4.210 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 3.840 1.790 4.000 ;
        RECT  1.630 3.840 1.790 4.460 ;
        RECT  1.630 4.300 2.020 4.460 ;
        RECT  0.660 3.840 0.860 4.490 ;
        RECT  0.580 2.810 2.060 2.970 ;
        RECT  0.140 1.450 2.680 1.610 ;
        RECT  0.140 1.450 0.340 1.810 ;
        RECT  0.140 0.300 1.530 0.460 ;
        RECT  1.370 0.300 1.530 0.640 ;
        RECT  1.370 0.480 3.220 0.640 ;
        RECT  0.140 0.300 0.340 0.650 ;
        RECT  0.660 0.620 0.940 0.960 ;
        RECT  0.660 0.800 3.790 0.960 ;
        RECT  3.630 0.800 3.790 1.620 ;
        RECT  2.950 1.460 3.790 1.620 ;
        RECT  2.950 1.460 3.110 1.990 ;
        RECT  0.580 1.770 3.110 1.990 ;
        RECT  2.250 2.810 3.170 2.970 ;
        RECT  3.010 2.810 3.170 3.300 ;
        RECT  3.010 3.140 3.970 3.300 ;
        RECT  3.810 3.140 3.970 4.000 ;
        RECT  3.150 3.840 3.970 4.000 ;
        RECT  3.150 3.840 3.310 4.460 ;
        RECT  2.250 4.300 3.310 4.460 ;
        LAYER VTPH ;
        RECT  2.080 1.090 2.880 3.660 ;
        RECT  0.000 1.140 4.400 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 4.400 4.800 ;
        RECT  0.000 0.000 4.400 1.090 ;
        RECT  0.000 0.000 2.080 1.140 ;
        RECT  2.880 0.000 4.400 1.140 ;
    END
END ADFM2HM

MACRO ADFM1HM
    CLASS CORE ;
    FOREIGN ADFM1HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.299  LAYER ME1  ;
        ANTENNADIFFAREA 0.299  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.010 4.200 4.210 4.400 ;
        LAYER ME2 ;
        RECT  3.910 4.000 4.300 4.400 ;
        LAYER ME1 ;
        RECT  3.910 4.200 4.300 4.500 ;
        RECT  4.130 2.820 4.300 4.500 ;
        RECT  3.970 2.820 4.300 3.030 ;
        END
    END S
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 3.400 1.280 ;
        RECT  0.100 0.840 0.360 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.374  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.830 3.520 3.590 3.680 ;
        RECT  2.010 3.980 2.990 4.140 ;
        RECT  2.830 3.520 2.990 4.140 ;
        RECT  2.010 3.460 2.300 4.140 ;
        RECT  1.340 3.460 2.300 3.640 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.281  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.490 3.130 2.650 3.780 ;
        RECT  0.480 3.130 2.650 3.290 ;
        RECT  0.480 3.130 0.700 3.680 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.296  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.980 0.390 4.300 1.750 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.450 2.260 3.730 2.970 ;
        RECT  3.350 1.780 3.630 2.540 ;
        RECT  0.140 2.260 0.340 3.030 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.460 -0.140 3.660 0.640 ;
        RECT  1.750 -0.140 2.030 0.320 ;
        RECT  0.000 4.660 4.400 4.940 ;
        RECT  3.490 4.240 3.690 4.940 ;
        RECT  1.180 4.220 1.380 4.940 ;
        RECT  0.140 4.210 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 3.840 1.790 4.000 ;
        RECT  1.630 3.840 1.790 4.460 ;
        RECT  1.630 4.300 2.020 4.460 ;
        RECT  0.660 3.840 0.860 4.490 ;
        RECT  0.580 2.810 2.060 2.970 ;
        RECT  0.140 1.450 2.680 1.610 ;
        RECT  0.140 1.450 0.340 1.980 ;
        RECT  0.140 0.300 1.530 0.460 ;
        RECT  1.370 0.300 1.530 0.640 ;
        RECT  1.370 0.480 3.220 0.640 ;
        RECT  0.140 0.300 0.340 0.650 ;
        RECT  0.660 0.620 0.940 0.960 ;
        RECT  0.660 0.800 3.790 0.960 ;
        RECT  3.630 0.800 3.790 1.620 ;
        RECT  2.950 1.460 3.790 1.620 ;
        RECT  2.950 1.460 3.110 1.990 ;
        RECT  0.580 1.770 3.110 1.990 ;
        RECT  2.250 2.810 3.170 2.970 ;
        RECT  3.010 2.810 3.170 3.360 ;
        RECT  3.010 3.200 3.970 3.360 ;
        RECT  3.810 3.200 3.970 4.000 ;
        RECT  3.150 3.840 3.970 4.000 ;
        RECT  3.150 3.840 3.310 4.460 ;
        RECT  2.250 4.300 3.310 4.460 ;
        LAYER VTPH ;
        RECT  2.080 1.090 2.880 3.660 ;
        RECT  0.000 1.140 4.400 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 4.400 4.800 ;
        RECT  0.000 0.000 4.400 1.090 ;
        RECT  0.000 0.000 2.080 1.140 ;
        RECT  2.880 0.000 4.400 1.140 ;
    END
END ADFM1HM

MACRO ADFM0HM
    CLASS CORE ;
    FOREIGN ADFM0HM 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 4.800 ;
    SYMMETRY X Y ;
    SITE CORE_6T2 ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        ANTENNADIFFAREA 0.235  LAYER ME2  ;
        PORT
        LAYER VI1 ;
        RECT  4.010 4.200 4.210 4.400 ;
        LAYER ME2 ;
        RECT  3.910 4.000 4.300 4.400 ;
        LAYER ME1 ;
        RECT  3.910 4.200 4.300 4.500 ;
        RECT  4.130 2.820 4.300 4.500 ;
        RECT  3.970 2.820 4.300 3.030 ;
        END
    END S
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.360  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  0.100 1.120 3.400 1.280 ;
        RECT  0.100 0.840 0.360 1.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.360  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.830 3.520 3.590 3.680 ;
        RECT  2.010 3.980 2.990 4.140 ;
        RECT  2.830 3.520 2.990 4.140 ;
        RECT  2.010 3.460 2.300 4.140 ;
        RECT  1.340 3.460 2.300 3.640 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  2.490 3.130 2.650 3.780 ;
        RECT  0.480 3.130 2.650 3.290 ;
        RECT  0.480 3.130 0.700 3.680 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.235  LAYER ME1  ;
        PORT
        LAYER ME1 ;
        RECT  3.980 0.390 4.300 1.750 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 2.260 4.400 2.540 ;
        RECT  3.450 2.260 3.730 2.970 ;
        RECT  3.350 1.780 3.630 2.540 ;
        RECT  0.140 2.260 0.340 3.030 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER ME1 ;
        RECT  0.000 -0.140 4.400 0.140 ;
        RECT  3.420 -0.140 3.700 0.640 ;
        RECT  1.750 -0.140 2.030 0.320 ;
        RECT  0.000 4.660 4.400 4.940 ;
        RECT  3.490 4.240 3.690 4.940 ;
        RECT  1.180 4.220 1.380 4.940 ;
        RECT  0.140 4.210 0.340 4.940 ;
        END
    END VSS
    OBS
        LAYER ME1 ;
        RECT  0.660 3.840 1.790 4.000 ;
        RECT  1.630 3.840 1.790 4.460 ;
        RECT  1.630 4.300 2.020 4.460 ;
        RECT  0.660 3.840 0.860 4.490 ;
        RECT  0.580 2.810 2.060 2.970 ;
        RECT  0.140 1.450 2.680 1.610 ;
        RECT  0.140 1.450 0.340 1.980 ;
        RECT  0.140 0.300 1.530 0.460 ;
        RECT  1.370 0.300 1.530 0.640 ;
        RECT  1.370 0.480 3.220 0.640 ;
        RECT  0.140 0.300 0.340 0.670 ;
        RECT  0.660 0.620 0.940 0.960 ;
        RECT  0.660 0.800 3.790 0.960 ;
        RECT  3.630 0.800 3.790 1.620 ;
        RECT  2.950 1.460 3.790 1.620 ;
        RECT  2.950 1.460 3.110 1.990 ;
        RECT  0.580 1.770 3.110 1.990 ;
        RECT  2.250 2.810 3.170 2.970 ;
        RECT  3.010 2.810 3.170 3.360 ;
        RECT  3.010 3.200 3.970 3.360 ;
        RECT  3.810 3.200 3.970 4.000 ;
        RECT  3.150 3.840 3.970 4.000 ;
        RECT  3.150 3.840 3.310 4.460 ;
        RECT  2.250 4.300 3.310 4.460 ;
        LAYER VTPH ;
        RECT  2.080 1.090 2.880 3.660 ;
        RECT  0.000 1.140 4.400 3.660 ;
        LAYER VTNH ;
        RECT  0.000 3.660 4.400 4.800 ;
        RECT  0.000 0.000 4.400 1.090 ;
        RECT  0.000 0.000 2.080 1.140 ;
        RECT  2.880 0.000 4.400 1.140 ;
    END
END ADFM0HM

END LIBRARY
