                                                           
.subckt ADFM0HM CO S A B CI VDD VSS 
MN0 net090 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net090 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net21 CI net090 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net21 A net084 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net084 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net096 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 net096 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net096 CI VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 net093 net21 net096 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN9 net0108 A net0111 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN10 net0111 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN11 net093 CI net0108 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 S net093 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN13 CO net21 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A net048 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD B net048 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net048 CI net21 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 net052 A net21 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B net052 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD A net054 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 VDD B net054 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD CI net054 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP8 net054 net21 net093 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP9 net064 A net067 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP10 VDD B net064 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP11 net067 CI net093 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP12 VDD net093 S VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP13 VDD net21 CO VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends ADFM0HM
                                                           
.subckt ADFM1HM CO S A B CI VDD VSS 
MN0 net090 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net090 B VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN2 net21 CI net090 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN3 net21 A net084 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN4 net084 B VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN5 net096 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 net096 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net096 CI VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 net093 net21 net096 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN9 net0108 A net0111 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN10 net0111 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN11 net093 CI net0108 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 S net093 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN13 CO net21 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net048 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 VDD B net048 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net048 CI net21 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 net052 A net21 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 VDD B net052 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP5 VDD A net054 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 VDD B net054 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD CI net054 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP8 net054 net21 net093 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP9 net064 A net067 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP10 VDD B net064 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP11 net067 CI net093 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP12 VDD net093 S VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP13 VDD net21 CO VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends ADFM1HM
                                                           
.subckt ADFM2HM CO S A B CI VDD VSS 
MN0 net090 A VSS VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN1 net090 B VSS VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN2 net21 CI net090 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN3 net21 A net084 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN4 net084 B VSS VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN5 net096 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 net096 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net096 CI VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 net093 net21 net096 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN9 net0108 A net0111 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN10 net0111 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN11 net093 CI net0108 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 S net093 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 CO net21 VSS VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MP0 VDD A net048 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP1 VDD B net048 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 net048 CI net21 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP3 net052 A net21 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP4 VDD B net052 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP5 VDD A net054 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD B net054 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP7 VDD CI net054 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP8 net054 net21 net093 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP9 net064 A net067 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP10 VDD B net064 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP11 net067 CI net093 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP12 VDD net093 S VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 VDD net21 CO VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends ADFM2HM
                                                           
.subckt ADFM4HM CO S A B CI VDD VSS 
MN0 net090 A VSS VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN1 net090 B VSS VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN2 net21 CI net090 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net21 A net084 VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN4 net084 B VSS VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN5 net096 A VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN6 net096 B VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net096 CI VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN8 net093 net21 net096 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0108 A net0111 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN10 net0111 B VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN11 net093 CI net0108 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN12 S net093 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 CO net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net048 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP1 VDD B net048 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net048 CI net21 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net052 A net21 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD B net052 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD A net054 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP6 VDD B net054 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP7 VDD CI net054 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP8 net054 net21 net093 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP9 net064 A net067 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP10 VDD B net064 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP11 net067 CI net093 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP12 VDD net093 S VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 VDD net21 CO VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends ADFM4HM
                                                           
.subckt ADFM8HM CO S A B CI VDD VSS 
MN0 net090 A VSS VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN1 net090 B VSS VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN2 net21 CI net090 VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN3 net21 A net084 VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN4 net084 B VSS VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN5 net096 A VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN6 net096 B VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN7 net096 CI VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN8 net093 net21 net096 VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN9 net0108 A net0111 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net0111 B VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN11 net093 CI net0108 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN12 S net093 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN13 CO net21 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A net048 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net048 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP2 net048 CI net21 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net052 A net21 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B net052 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD A net054 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP6 VDD B net054 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP7 VDD CI net054 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP8 net054 net21 net093 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP9 net064 A net067 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD B net064 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net067 CI net093 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net093 S VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 VDD net21 CO VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends ADFM8HM
                                                           
.subckt ADHM0HM CO S A B VDD VSS 
MN0 net01 A net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net05 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 net01 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 S net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 CO net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 net04 A net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net03 S VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP6 VDD net01 CO VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends ADHM0HM
                                                           
.subckt ADHM1HM CO S A B VDD VSS 
MN0 net01 A net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net05 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 net01 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 S net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN6 CO net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.30u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.30u l=0.12u
MP2 net04 A net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net03 S VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP6 VDD net01 CO VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends ADHM1HM
                                                           
.subckt ADHM2HM CO S A B VDD VSS 
MN0 net01 A net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN2 net05 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 net01 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 S net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 CO net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP2 net04 A net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net03 S VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net01 CO VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends ADHM2HM
                                                           
.subckt ADHM4HM CO S A B VDD VSS 
MN0 net01 A net02 VSS N_15_LL_EE2_UCFN w=0.7u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.7u l=0.12u
MN2 net05 A VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net03 net01 net05 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN5 S net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN6 CO net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP2 net04 A net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP5 VDD net03 S VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net01 CO VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends ADHM4HM
                                                           
.subckt ADHM8HM CO S A B VDD VSS 
MN0 net01 A net02 VSS N_15_LL_EE2_UCFN w=0.72u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.72u l=0.12u
MN2 net05 A VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN4 net03 net01 net05 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN5 S net03 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN6 CO net01 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP2 net04 A net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD net03 S VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP6 VDD net01 CO VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends ADHM8HM
                                                           
.subckt AN2M0HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AN2M0HM
                                                           
.subckt AN2M12HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends AN2M12HM
                                                           
.subckt AN2M16HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=1.81u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.81u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends AN2M16HM
                                                           
.subckt AN2M1HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AN2M1HM
                                                           
.subckt AN2M2HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AN2M2HM
                                                           
.subckt AN2M4HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AN2M4HM
                                                           
.subckt AN2M6HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends AN2M6HM
                                                           
.subckt AN2M8HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=1.03u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.03u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AN2M8HM
                                                           
.subckt AN3M0HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AN3M0HM
                                                           
.subckt AN3M12HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends AN3M12HM
                                                           
.subckt AN3M16HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends AN3M16HM
                                                           
.subckt AN3M1HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AN3M1HM
                                                           
.subckt AN3M2HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AN3M2HM
                                                           
.subckt AN3M4HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AN3M4HM
                                                           
.subckt AN3M6HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends AN3M6HM
                                                           
.subckt AN3M8HM Z A B C VDD VSS 
MN0 net03 A net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 B net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A net03 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP1 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AN3M8HM
                                                           
.subckt AN4M0HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AN4M0HM
                                                           
.subckt AN4M12HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends AN4M12HM
                                                           
.subckt AN4M16HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=1.98u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=1.57u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends AN4M16HM
                                                           
.subckt AN4M1HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AN4M1HM
                                                           
.subckt AN4M2HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AN4M2HM
                                                           
.subckt AN4M4HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AN4M4HM
                                                           
.subckt AN4M6HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends AN4M6HM
                                                           
.subckt AN4M8HM Z A B C D VDD VSS 
MN0 net04 A net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 B net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 C net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net04 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP4 VDD net04 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AN4M8HM
                                                           
.subckt ANTHM A VDD VSS 
DZ0 VSS A DION_EE2_UCFN area=0.372p pj=2.44u
.ends ANTHM
                                                           
.subckt AO211M0HM Z A1 A2 B C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO211M0HM
                                                           
.subckt AO211M1HM Z A1 A2 B C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO211M1HM
                                                           
.subckt AO211M2HM Z A1 A2 B C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO211M2HM
                                                           
.subckt AO211M4HM Z A1 A2 B C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO211M4HM
                                                           
.subckt AO211M8HM Z A1 A2 B C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO211M8HM
                                                           
.subckt AO21M0HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO21M0HM
                                                           
.subckt AO21M1HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO21M1HM
                                                           
.subckt AO21M2HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO21M2HM
                                                           
.subckt AO21M4HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO21M4HM
                                                           
.subckt AO21M8HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=1.03u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=1.03u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO21M8HM
                                                           
.subckt AO221M0HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO221M0HM
                                                           
.subckt AO221M1HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO221M1HM
                                                           
.subckt AO221M2HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO221M2HM
                                                           
.subckt AO221M4HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO221M4HM
                                                           
.subckt AO221M8HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO221M8HM
                                                           
.subckt AO222M0HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD C1 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD C2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO222M0HM
                                                           
.subckt AO222M1HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD C1 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD C2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO222M1HM
                                                           
.subckt AO222M2HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD C1 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD C2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO222M2HM
                                                           
.subckt AO222M4HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net01 C1 net06 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net06 C2 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD C2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO222M4HM
                                                           
.subckt AO222M8HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net01 A1 net04 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 net04 A2 VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN2 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN3 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN4 net01 C1 net06 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN5 net06 C2 VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP2 net03 B1 net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP3 net03 B2 net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP4 VDD C1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD C2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO222M8HM
                                                           
.subckt AO22B10M0HM Z A1 B1 B2 NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net03 net01 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO22B10M0HM
                                                           
.subckt AO22B10M1HM Z A1 B1 B2 NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net03 net01 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO22B10M1HM
                                                           
.subckt AO22B10M2HM Z A1 B1 B2 NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net03 net01 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO22B10M2HM
                                                           
.subckt AO22B10M4HM Z A1 B1 B2 NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A1 net04 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net02 B1 net05 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 net01 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO22B10M4HM
                                                           
.subckt AO22B10M8HM Z A1 B1 B2 NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN1 net02 A1 net04 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 net02 B1 net05 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net03 net01 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO22B10M8HM
                                                           
.subckt AO22B11M0HM Z A1 B1 NA2 NB2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 NB2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 A1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 B1 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD NB2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B1 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO22B11M0HM
                                                           
.subckt AO22B11M1HM Z A1 B1 NA2 NB2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 NB2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 A1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 B1 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD NB2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B1 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO22B11M1HM
                                                           
.subckt AO22B11M2HM Z A1 B1 NA2 NB2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 NB2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 A1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 B1 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD NB2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B1 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO22B11M2HM
                                                           
.subckt AO22B11M4HM Z A1 B1 NA2 NB2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 NB2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net05 A1 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net03 net01 net05 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net06 B1 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN5 net03 net02 net06 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD NB2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B1 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net02 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO22B11M4HM
                                                           
.subckt AO22B11M8HM Z A1 B1 NA2 NB2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN1 net02 NB2 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN2 net03 A1 net05 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 net03 B1 net06 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN5 net06 net02 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 VDD NB2 net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD B1 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD net02 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO22B11M8HM
                                                           
.subckt AO22M0HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO22M0HM
                                                           
.subckt AO22M1HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO22M1HM
                                                           
.subckt AO22M2HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO22M2HM
                                                           
.subckt AO22M4HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net01 B1 net04 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO22M4HM
                                                           
.subckt AO22M8HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN2 net01 B1 net04 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO22M8HM
                                                           
.subckt AO31M0HM Z A1 A2 A3 B VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO31M0HM
                                                           
.subckt AO31M1HM Z A1 A2 A3 B VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO31M1HM
                                                           
.subckt AO31M2HM Z A1 A2 A3 B VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO31M2HM
                                                           
.subckt AO31M4HM Z A1 A2 A3 B VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO31M4HM
                                                           
.subckt AO31M8HM Z A1 A2 A3 B VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO31M8HM
                                                           
.subckt AO32M0HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO32M0HM
                                                           
.subckt AO32M1HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO32M1HM
                                                           
.subckt AO32M2HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO32M2HM
                                                           
.subckt AO32M4HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO32M4HM
                                                           
.subckt AO32M8HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 net05 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO32M8HM
                                                           
.subckt AO33M0HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD B3 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AO33M0HM
                                                           
.subckt AO33M1HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD B3 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AO33M1HM
                                                           
.subckt AO33M2HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 B2 net06 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net06 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD B3 net02 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AO33M2HM
                                                           
.subckt AO33M4HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net05 B2 net06 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net06 B3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD B3 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AO33M4HM
                                                           
.subckt AO33M8HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net01 A1 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 A2 net04 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net04 A3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 B1 net05 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net05 B2 net06 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net06 B3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN6 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net02 A2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 A3 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD B3 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AO33M8HM
                                                           
.subckt AOI211M0HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 Z C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI211M0HM
                                                           
.subckt AOI211M1HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN3 Z C VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP2 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP3 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
.ends AOI211M1HM
                                                           
.subckt AOI211M2HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 Z C VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI211M2HM
                                                           
.subckt AOI211M4HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.88u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.88u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 B net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD C net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI211M4HM
                                                           
.subckt AOI211M8HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.76u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=1.76u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 Z C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net02 B net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD C net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI211M8HM
                                                           
.subckt AOI21B01M0HM Z A1 A2 NB VDD VSS 
MN0 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP0 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net02 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI21B01M0HM
                                                           
.subckt AOI21B01M1HM Z A1 A2 NB VDD VSS 
MN0 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net02 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI21B01M1HM
                                                           
.subckt AOI21B01M2HM Z A1 A2 NB VDD VSS 
MN0 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI21B01M2HM
                                                           
.subckt AOI21B01M4HM Z A1 A2 NB VDD VSS 
MN0 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN2 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MP0 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI21B01M4HM
                                                           
.subckt AOI21B01M8HM Z A1 A2 NB VDD VSS 
MN0 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.89u l=0.12u
MN2 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=1.89u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.32u l=0.12u
MP0 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net02 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI21B01M8HM
                                                           
.subckt AOI21B10M0HM Z A1 B NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net02 net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI21B10M0HM
                                                           
.subckt AOI21B10M1HM Z A1 B NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net02 net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI21B10M1HM
                                                           
.subckt AOI21B10M2HM Z A1 B NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI21B10M2HM
                                                           
.subckt AOI21B10M4HM Z A1 B NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN2 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI21B10M4HM
                                                           
.subckt AOI21B10M8HM Z A1 B NA2 VDD VSS 
MN0 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.89u l=0.12u
MN2 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=1.89u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=1.32u l=0.12u
MP0 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net02 net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI21B10M8HM
                                                           
.subckt AOI21B20M0HM Z B NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net03 B Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI21B20M0HM
                                                           
.subckt AOI21B20M1HM Z B NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net03 B Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI21B20M1HM
                                                           
.subckt AOI21B20M2HM Z B NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI21B20M2HM
                                                           
.subckt AOI21B20M4HM Z B NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net03 B Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI21B20M4HM
                                                           
.subckt AOI21B20M8HM Z B NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net03 B Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI21B20M8HM
                                                           
.subckt AOI21M0HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI21M0HM
                                                           
.subckt AOI21M1HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI21M1HM
                                                           
.subckt AOI21M2HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI21M2HM
                                                           
.subckt AOI21M3HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.80u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.80u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
.ends AOI21M3HM
                                                           
.subckt AOI21M4HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI21M4HM
                                                           
.subckt AOI21M6HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends AOI21M6HM
                                                           
.subckt AOI21M8HM Z A1 A2 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN2 Z B VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD B net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI21M8HM
                                                           
.subckt AOI221M0HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN4 Z C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI221M0HM
                                                           
.subckt AOI221M1HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z C VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI221M1HM
                                                           
.subckt AOI221M2HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 Z C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI221M2HM
                                                           
.subckt AOI221M4HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN4 Z C VSS VSS N_15_LL_EE2_UCFN w=0.63u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD C net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI221M4HM
                                                           
.subckt AOI221M8HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN4 Z C VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD C net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI221M8HM
                                                           
.subckt AOI222M0HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN4 Z C1 net05 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN5 net05 C2 VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD C1 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 VDD C2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI222M0HM
                                                           
.subckt AOI222M1HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z C1 net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net05 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD C1 net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD C2 net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI222M1HM
                                                           
.subckt AOI222M2HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 Z C1 net05 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net05 C2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD C2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI222M2HM
                                                           
.subckt AOI222M4HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN4 Z C1 net05 VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MN5 net05 C2 VSS VSS N_15_LL_EE2_UCFN w=0.87u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD C1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD C2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI222M4HM
                                                           
.subckt AOI222M8HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN1 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN2 Z B1 net04 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN4 Z C1 net05 VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MN5 net05 C2 VSS VSS N_15_LL_EE2_UCFN w=1.75u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net02 B2 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD C1 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 VDD C2 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI222M8HM
                                                           
.subckt AOI22B20M0HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net03 B2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net03 B1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI22B20M0HM
                                                           
.subckt AOI22B20M1HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net03 B2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 net03 B1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI22B20M1HM
                                                           
.subckt AOI22B20M2HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net03 B2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net03 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI22B20M2HM
                                                           
.subckt AOI22B20M4HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net03 B2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net03 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI22B20M4HM
                                                           
.subckt AOI22B20M8HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net01 NA1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net02 NA1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net03 B2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 net03 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI22B20M8HM
                                                           
.subckt AOI22M0HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net03 B2 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI22M0HM
                                                           
.subckt AOI22M1HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net03 B2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
.ends AOI22M1HM
                                                           
.subckt AOI22M2HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net03 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI22M2HM
                                                           
.subckt AOI22M4HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 net03 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI22M4HM
                                                           
.subckt AOI22M8HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN3 net03 B2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI22M8HM
                                                           
.subckt AOI31M0HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI31M0HM
                                                           
.subckt AOI31M1HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI31M1HM
                                                           
.subckt AOI31M2HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI31M2HM
                                                           
.subckt AOI31M4HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI31M4HM
                                                           
.subckt AOI31M8HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MN3 Z B VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI31M8HM
                                                           
.subckt AOI32M0HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI32M0HM
                                                           
.subckt AOI32M1HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI32M1HM
                                                           
.subckt AOI32M2HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI32M2HM
                                                           
.subckt AOI32M4HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI32M4HM
                                                           
.subckt AOI32M8HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN4 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI32M8HM
                                                           
.subckt AOI33M0HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net04 B2 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN5 net05 B3 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 VDD B3 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends AOI33M0HM
                                                           
.subckt AOI33M1HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN4 net04 B2 net05 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN5 net05 B3 VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD B3 net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends AOI33M1HM
                                                           
.subckt AOI33M2HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net04 B2 net05 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net05 B3 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD B3 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends AOI33M2HM
                                                           
.subckt AOI33M4HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net04 B2 net05 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net05 B3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD B3 net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends AOI33M4HM
                                                           
.subckt AOI33M8HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 net02 A2 net03 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net03 A3 VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MN3 Z B1 net04 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN4 net04 B2 net05 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN5 net05 B3 VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MP0 net01 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net01 A2 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net01 A3 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 VDD B3 net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends AOI33M8HM
                                                           
.subckt BHDM1HM Z VDD VSS 
MN0 net9 Z VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN1 Z net9 net3 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net3 net9 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD Z net9 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP1 VDD net9 Z VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends BHDM1HM
                                                           
.subckt BUFM10HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.80u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.15u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=3.40u l=0.12u
.ends BUFM10HM
                                                           
.subckt BUFM12HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends BUFM12HM
                                                           
.subckt BUFM14HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=3.92u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=4.76u l=0.12u
.ends BUFM14HM
                                                           
.subckt BUFM16HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends BUFM16HM
                                                           
.subckt BUFM18HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=5.04u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=6.12u l=0.12u
.ends BUFM18HM
                                                           
.subckt BUFM20HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=5.60u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=6.80u l=0.12u
.ends BUFM20HM
                                                           
.subckt BUFM24HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=6.72u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
.ends BUFM24HM
                                                           
.subckt BUFM28HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=7.84u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=9.52u l=0.12u
.ends BUFM28HM
                                                           
.subckt BUFM2HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends BUFM2HM
                                                           
.subckt BUFM32HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=8.96u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
.ends BUFM32HM
                                                           
.subckt BUFM36HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=2.80u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=10.08u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=3.40u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=12.24u l=0.12u
.ends BUFM36HM
                                                           
.subckt BUFM3HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
.ends BUFM3HM
                                                           
.subckt BUFM40HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=2.80u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=10.64u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=3.40u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=12.92u l=0.12u
.ends BUFM40HM
                                                           
.subckt BUFM48HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=12.88u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=15.64u l=0.12u
.ends BUFM48HM
                                                           
.subckt BUFM4HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends BUFM4HM
                                                           
.subckt BUFM5HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.41u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.72u l=0.12u
.ends BUFM5HM
                                                           
.subckt BUFM6HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends BUFM6HM
                                                           
.subckt BUFM8HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends BUFM8HM
                                                           
.subckt BUFTM12HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends BUFTM12HM
                                                           
.subckt BUFTM16HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=1.36u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.68u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=1.68u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.86u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=5.42u l=0.12u
.ends BUFTM16HM
                                                           
.subckt BUFTM1HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends BUFTM1HM
                                                           
.subckt BUFTM20HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.63u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=1.88u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=5.60u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.76u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=2.29u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=1.15u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=6.80u l=0.12u
.ends BUFTM20HM
                                                           
.subckt BUFTM24HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=6.24u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=8u l=0.12u
.ends BUFTM24HM
                                                           
.subckt BUFTM2HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends BUFTM2HM
                                                           
.subckt BUFTM3HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
.ends BUFTM3HM
                                                           
.subckt BUFTM4HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends BUFTM4HM
                                                           
.subckt BUFTM6HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends BUFTM6HM
                                                           
.subckt BUFTM8HM Z A E VDD VSS 
MN0 net36 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net45 net36 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net45 A VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN3 net45 E net55 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN4 Z net45 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD E net36 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD E net55 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A net55 VDD P_15_LL_EE2_UCFN w=0.89u l=0.12u
MP3 net55 net36 net45 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP4 VDD net55 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends BUFTM8HM
                                                           
.subckt CKAN2M12HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends CKAN2M12HM
                                                           
.subckt CKAN2M16HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.61u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=1.4u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.4u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends CKAN2M16HM
                                                           
.subckt CKAN2M2HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKAN2M2HM
                                                           
.subckt CKAN2M3HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.05u l=0.12u
.ends CKAN2M3HM
                                                           
.subckt CKAN2M4HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.65u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends CKAN2M4HM
                                                           
.subckt CKAN2M6HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends CKAN2M6HM
                                                           
.subckt CKAN2M8HM Z A B VDD VSS 
MN0 net02 A net01 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN2 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.31u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends CKAN2M8HM
                                                           
.subckt CKBUFM12HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.57u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.7u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends CKBUFM12HM
                                                           
.subckt CKBUFM16HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.76u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.27u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.82u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends CKBUFM16HM
                                                           
.subckt CKBUFM1HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends CKBUFM1HM
                                                           
.subckt CKBUFM20HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.83u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.26u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=6.8u l=0.12u
.ends CKBUFM20HM
                                                           
.subckt CKBUFM24HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.13u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=3.4u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
.ends CKBUFM24HM
                                                           
.subckt CKBUFM2HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKBUFM2HM
                                                           
.subckt CKBUFM32HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.5u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=4.53u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=3.62u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
.ends CKBUFM32HM
                                                           
.subckt CKBUFM3HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
.ends CKBUFM3HM
                                                           
.subckt CKBUFM40HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.9u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=5.67u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=4.54u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=13.6u l=0.12u
.ends CKBUFM40HM
                                                           
.subckt CKBUFM48HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=2.26u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=6.8u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=16.32u l=0.12u
.ends CKBUFM48HM
                                                           
.subckt CKBUFM4HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends CKBUFM4HM
                                                           
.subckt CKBUFM6HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends CKBUFM6HM
                                                           
.subckt CKBUFM8HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN1 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.14u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP1 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends CKBUFM8HM
                                                           
.subckt CKINVM12HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.7u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends CKINVM12HM
                                                           
.subckt CKINVM16HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.26u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends CKINVM16HM
                                                           
.subckt CKINVM1HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends CKINVM1HM
                                                           
.subckt CKINVM20HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.83u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=6.8u l=0.12u
.ends CKINVM20HM
                                                           
.subckt CKINVM24HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=3.4u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
.ends CKINVM24HM
                                                           
.subckt CKINVM2HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKINVM2HM
                                                           
.subckt CKINVM32HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=4.53u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
.ends CKINVM32HM
                                                           
.subckt CKINVM3HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
.ends CKINVM3HM
                                                           
.subckt CKINVM40HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=5.67u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=13.6u l=0.12u
.ends CKINVM40HM
                                                           
.subckt CKINVM48HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=6.8u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=16.32u l=0.12u
.ends CKINVM48HM
                                                           
.subckt CKINVM4HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.57u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends CKINVM4HM
                                                           
.subckt CKINVM6HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends CKINVM6HM
                                                           
.subckt CKINVM8HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.13u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends CKINVM8HM
                                                           
.subckt CKMUX2M12HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=1.74u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
.ends CKMUX2M12HM
                                                           
.subckt CKMUX2M2HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
.ends CKMUX2M2HM
                                                           
.subckt CKMUX2M3HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKMUX2M3HM
                                                           
.subckt CKMUX2M4HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=0.65u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKMUX2M4HM
                                                           
.subckt CKMUX2M6HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=0.97u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKMUX2M6HM
                                                           
.subckt CKMUX2M8HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=1.30u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKMUX2M8HM
                                                           
.subckt CKND2M12HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=2.5u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=2.5u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends CKND2M12HM
                                                           
.subckt CKND2M16HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=3.94u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=3.94u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends CKND2M16HM
                                                           
.subckt CKND2M2HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends CKND2M2HM
                                                           
.subckt CKND2M4HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends CKND2M4HM
                                                           
.subckt CKND2M6HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends CKND2M6HM
                                                           
.subckt CKND2M8HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.97u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.97u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends CKND2M8HM
                                                           
.subckt CKXOR2M12HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.88u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=1.7u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=1.08u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=1.06u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=1.06u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends CKXOR2M12HM
                                                           
.subckt CKXOR2M1HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends CKXOR2M1HM
                                                           
.subckt CKXOR2M2HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
.ends CKXOR2M2HM
                                                           
.subckt CKXOR2M4HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends CKXOR2M4HM
                                                           
.subckt CKXOR2M8HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.64u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=1.17u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.26u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=2.68u l=0.12u
.ends CKXOR2M8HM
                                                           
.subckt DEL1M1HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends DEL1M1HM
                                                           
.subckt DEL1M4HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends DEL1M4HM
                                                           
.subckt DEL2M1HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.24u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.24u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.22u l=0.24u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.22u l=0.24u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends DEL2M1HM
                                                           
.subckt DEL2M4HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.24u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.24u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.47u l=0.24u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.47u l=0.24u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends DEL2M4HM
                                                           
.subckt DEL3M1HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.36u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.36u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.22u l=0.36u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.22u l=0.36u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends DEL3M1HM
                                                           
.subckt DEL3M4HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.36u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.36u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.47u l=0.36u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.47u l=0.36u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends DEL3M4HM
                                                           
.subckt DEL4M1HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.48u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.48u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.22u l=0.48u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.22u l=0.48u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends DEL4M1HM
                                                           
.subckt DEL4M4HM Z A VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.48u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.48u
MN3 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP1 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.47u l=0.48u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.47u l=0.48u
MP3 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends DEL4M4HM
                                                           
.subckt DFCM1HM Q QB CKB D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFCM1HM
                                                           
.subckt DFCM2HM Q QB CKB D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFCM2HM
                                                           
.subckt DFCM4HM Q QB CKB D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFCM4HM
                                                           
.subckt DFCM8HM Q QB CKB D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFCM8HM
                                                           
.subckt DFCQM1HM Q CKB D VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFCQM1HM
                                                           
.subckt DFCQM2HM Q CKB D VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFCQM2HM
                                                           
.subckt DFCQM4HM Q CKB D VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFCQM4HM
                                                           
.subckt DFCQM8HM Q CKB D VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFCQM8HM
                                                           
.subckt DFCQRSM1HM Q CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.43u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.43u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFCQRSM1HM
                                                           
.subckt DFCQRSM2HM Q CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFCQRSM2HM
                                                           
.subckt DFCQRSM4HM Q CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFCQRSM4HM
                                                           
.subckt DFCQRSM8HM Q CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.7u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.91u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFCQRSM8HM
                                                           
.subckt DFCRSM1HM Q QB CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.43u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.43u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFCRSM1HM
                                                           
.subckt DFCRSM2HM Q QB CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFCRSM2HM
                                                           
.subckt DFCRSM4HM Q QB CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFCRSM4HM
                                                           
.subckt DFCRSM8HM Q QB CKB D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.7u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP2 VDD CKB net11 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.91u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.91u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN1 net11 CKB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFCRSM8HM
                                                           
.subckt DFEM1HM Q QB CK D E VDD VSS 
MP22 net079 net0215 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net079 net0190 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 net0190 E net0187 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 net0187 net0130 net047 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP20 net0158 net0215 net0187 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP21 net019 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net11 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net0215 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 VDD D net047 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD CK net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net0128 net0215 net019 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN21 net0128 net11 net079 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net047 E net0244 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net0244 net0130 net0234 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net0234 net079 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net0244 net11 net0158 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0215 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0215 net11 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net047 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net11 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends DFEM1HM
                                                           
.subckt DFEM2HM Q QB CK D E VDD VSS 
MP22 net079 net0215 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net079 net0190 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP18 net0190 E net0187 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP19 net0187 net0130 net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP20 net0158 net0215 net0187 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net019 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net11 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net0215 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 VDD D net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD CK net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net0128 net0215 net019 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN21 net0128 net11 net079 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net047 E net0244 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN17 net0244 net0130 net0234 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN18 net0234 net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN19 net0244 net11 net0158 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0215 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0215 net11 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net047 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net11 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends DFEM2HM
                                                           
.subckt DFEM4HM Q QB CK D E VDD VSS 
MP22 net079 net0215 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net079 net0190 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP18 net0190 E net0187 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP19 net0187 net0130 net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP20 net0158 net0215 net0187 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net019 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net11 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net0215 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 VDD D net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD CK net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net0128 net0215 net019 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN21 net0128 net11 net079 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN16 net047 E net0244 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN17 net0244 net0130 net0234 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN18 net0234 net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN19 net0244 net11 net0158 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0215 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0215 net11 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net047 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN1 net11 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends DFEM4HM
                                                           
.subckt DFEM8HM Q QB CK D E VDD VSS 
MP22 net079 net0215 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net079 net0190 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP18 net0190 E net0187 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP19 net0187 net0130 net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP20 net0158 net0215 net0187 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net019 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net11 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net0215 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 VDD D net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD CK net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net0128 net0215 net019 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN21 net0128 net11 net079 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN16 net047 E net0244 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN17 net0244 net0130 net0234 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN18 net0234 net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN19 net0244 net11 net0158 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0215 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0215 net11 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net047 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN1 net11 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends DFEM8HM
                                                           
.subckt DFEQM1HM Q CK D E VDD VSS 
MN9 net0123 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0125 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net18 net0266 net13 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net15 net14 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net18 net0123 net15 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net0125 E net18 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net29 net13 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net13 net51 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net29 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net81 net51 net29 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net36 net81 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 Q net36 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN25 net81 net0266 net14 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net36 net14 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net51 net0266 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0266 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP8 VDD E net0123 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD D net0125 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net13 net51 net64 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net64 net0123 net0125 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net67 E net64 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 VDD net14 net67 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD net13 net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net79 net29 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net79 net0266 net13 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net29 net0266 net81 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net81 net36 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP19 VDD net36 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP29 net14 net36 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP26 net14 net51 net81 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0266 net51 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP4 VDD CK net0266 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
.ends DFEQM1HM
                                                           
.subckt DFEQM2HM Q CK D E VDD VSS 
MN9 net0123 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0125 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN6 net18 net0266 net13 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net15 net14 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net18 net0123 net15 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net0125 E net18 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN10 net29 net13 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net13 net51 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net29 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net81 net51 net29 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net36 net81 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN18 Q net36 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN25 net81 net0266 net14 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net36 net14 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net51 net0266 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0266 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP8 VDD E net0123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D net0125 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 net13 net51 net64 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net64 net0123 net0125 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net67 E net64 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 VDD net14 net67 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP12 VDD net13 net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net79 net29 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net79 net0266 net13 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net29 net0266 net81 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP16 VDD net81 net36 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD net36 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP29 net14 net36 VDD VDD P_15_LL_EE2_UCFN w=0.23u l=0.12u
MP26 net14 net51 net81 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0266 net51 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD CK net0266 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFEQM2HM
                                                           
.subckt DFEQM4HM Q CK D E VDD VSS 
MN9 net0123 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0125 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN6 net18 net0266 net13 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net15 net14 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net18 net0123 net15 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net0125 E net18 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN10 net29 net13 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net13 net51 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net29 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net81 net51 net29 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net36 net81 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN18 Q net36 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN25 net81 net0266 net14 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net36 net14 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net51 net0266 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0266 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP8 VDD E net0123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D net0125 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 net13 net51 net64 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net64 net0123 net0125 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net67 E net64 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD net14 net67 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP12 VDD net13 net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net79 net29 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net79 net0266 net13 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net29 net0266 net81 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP16 VDD net81 net36 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD net36 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP29 net14 net36 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net14 net51 net81 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0266 net51 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD CK net0266 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFEQM4HM
                                                           
.subckt DFEQM8HM Q CK D E VDD VSS 
MN9 net0123 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0125 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN6 net18 net0266 net13 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 net15 net14 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net18 net0123 net15 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net0125 E net18 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN10 net29 net13 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN12 net13 net51 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net29 net31 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net81 net51 net29 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN15 net36 net81 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN18 Q net36 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN25 net81 net0266 net14 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN29 VSS net36 net14 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net51 net0266 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0266 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP8 VDD E net0123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D net0125 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 net13 net51 net64 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net64 net0123 net0125 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net67 E net64 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD net14 net67 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP12 VDD net13 net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net79 net29 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net79 net0266 net13 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net29 net0266 net81 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP16 VDD net81 net36 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD net36 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP29 net14 net36 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net14 net51 net81 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0266 net51 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD CK net0266 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFEQM8HM
                                                           
.subckt DFEQRM1HM Q CK D E RB VDD VSS 
MN17 net42 net64 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net10 RB VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN16 net10 net12 net64 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN10 Q net64 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net42 net0295 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net29 net58 net25 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net25 net0295 net40 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net31 net27 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net31 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net12 net58 net27 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net0283 E net40 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net40 net0286 net43 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net43 net42 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0283 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net0286 E VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net27 net25 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net58 net0295 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0295 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP20 net27 net0295 net12 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP16 net64 net12 VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP15 VDD net64 net42 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP14 VDD net64 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP12 net12 net58 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net82 net27 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net82 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net42 net89 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net89 E net92 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net92 net0286 net0283 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net25 net58 net92 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D net0283 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP8 VDD E net0286 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD net25 net27 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP11 net82 net0295 net25 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0295 net58 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD CK net0295 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFEQRM1HM
                                                           
.subckt DFEQRM2HM Q CK D E RB VDD VSS 
MN17 net42 net64 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 net10 RB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN16 net10 net12 net64 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN10 Q net64 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN15 net42 net0295 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net29 net58 net25 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net25 net0295 net40 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN11 net31 net27 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net31 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net12 net58 net27 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0283 E net40 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net40 net0286 net43 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net43 net42 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net0283 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net0286 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net27 net25 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net58 net0295 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0295 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP20 net27 net0295 net12 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP16 net64 net12 VDD VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 VDD net64 net42 VDD P_15_LL_EE2_UCFN w=0.23u l=0.12u
MP14 VDD net64 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 net12 net58 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net82 net27 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net82 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net42 net89 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP3 net89 E net92 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP5 net92 net0286 net0283 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 net25 net58 net92 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP7 VDD D net0283 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD E net0286 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net25 net27 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP11 net82 net0295 net25 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0295 net58 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0295 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends DFEQRM2HM
                                                           
.subckt DFEQRM4HM Q CK D E RB VDD VSS 
MN17 net42 net64 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 net10 RB VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN16 net10 net12 net64 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN10 Q net64 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN15 net42 net0295 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net29 net58 net25 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net25 net0295 net40 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN11 net31 net27 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net31 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net12 net58 net27 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0283 E net40 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net40 net0286 net43 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net43 net42 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net0283 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net0286 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net27 net25 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net58 net0295 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0295 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP20 net27 net0295 net12 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 VDD RB net64 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP16 net64 net12 VDD VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP15 VDD net64 net42 VDD P_15_LL_EE2_UCFN w=0.23u l=0.12u
MP14 VDD net64 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP12 net12 net58 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net82 net27 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net82 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net42 net89 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP3 net89 E net92 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP5 net92 net0286 net0283 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 net25 net58 net92 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP7 VDD D net0283 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD E net0286 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net25 net27 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP11 net82 net0295 net25 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0295 net58 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0295 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends DFEQRM4HM
                                                           
.subckt DFEQRM8HM Q CK D E RB VDD VSS 
MN17 net42 net64 VSS VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN6 net10 RB VSS VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MN16 net10 net12 net64 VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MN10 Q net64 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN15 net42 net0295 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net29 net58 net25 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net25 net0295 net40 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN11 net31 net27 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net31 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net12 net58 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0283 E net40 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN3 net40 net0286 net43 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 net43 net42 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net0283 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN9 net0286 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net27 net25 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net58 net0295 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0295 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP20 net27 net0295 net12 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP17 VDD RB net64 VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP16 net64 net12 VDD VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP15 VDD net64 net42 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP14 VDD net64 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP12 net12 net58 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net82 net27 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP9 VDD RB net82 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD net42 net89 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net89 E net92 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net92 net0286 net0283 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 net25 net58 net92 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD D net0283 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD E net0286 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net25 net27 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net82 net0295 net25 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD net0295 net58 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP4 VDD CK net0295 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFEQRM8HM
                                                           
.subckt DFEQZRM1HM Q CK D E RB VDD VSS 
MP18 net20 net75 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD E net58 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP15 VDD RB net13 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP11 net13 net79 net61 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net20 E net13 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0301 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP1 VDD net0301 net79 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net61 net90 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net35 net90 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net35 net0301 net61 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net90 net0301 net37 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net37 net97 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD net97 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP29 net75 net97 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP26 net75 net79 net37 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net53 D net13 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD net58 net53 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MN16 net58 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN14 net61 net0301 net73 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN11 net71 RB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net73 net58 net77 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net70 E net71 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net73 D net70 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net71 net75 net77 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0301 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net79 net0301 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net90 net61 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net61 net79 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net90 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net37 net79 net90 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net97 net37 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 Q net97 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN25 net37 net0301 net75 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net97 net75 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends DFEQZRM1HM
                                                           
.subckt DFEQZRM2HM Q CK D E RB VDD VSS 
MP18 net20 net75 VDD VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP17 VDD E net58 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP15 VDD RB net13 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP11 net13 net79 net61 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net20 E net13 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP4 VDD CK net0301 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD net0301 net79 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net61 net90 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net35 net90 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net35 net0301 net61 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net90 net0301 net37 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP16 VDD net37 net97 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD net97 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP29 net75 net97 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net75 net79 net37 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net53 D net13 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD net58 net53 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MN16 net58 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 net61 net0301 net73 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN11 net71 RB VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net73 net58 net77 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net70 E net71 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net73 D net70 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN17 net71 net75 net77 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net0301 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net79 net0301 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net90 net61 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net61 net79 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net90 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net37 net79 net90 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net97 net37 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN18 Q net97 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN25 net37 net0301 net75 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net97 net75 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
.ends DFEQZRM2HM
                                                           
.subckt DFEQZRM4HM Q CK D E RB VDD VSS 
MP18 net20 net75 VDD VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP17 VDD E net58 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP15 VDD RB net13 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP11 net13 net79 net61 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net20 E net13 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP4 VDD CK net0301 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD net0301 net79 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net61 net90 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net35 net90 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net35 net0301 net61 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net90 net0301 net37 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP16 VDD net37 net97 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD net97 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP29 net75 net97 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net75 net79 net37 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net53 D net13 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD net58 net53 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MN16 net58 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 net61 net0301 net73 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN11 net71 RB VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net73 net58 net77 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net70 E net71 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net73 D net70 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN17 net71 net75 net77 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net0301 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net79 net0301 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net90 net61 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net61 net79 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net90 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net37 net79 net90 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net97 net37 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN18 Q net97 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN25 net37 net0301 net75 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net97 net75 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
.ends DFEQZRM4HM
                                                           
.subckt DFEQZRM8HM Q CK D E RB VDD VSS 
MP18 net20 net75 VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP17 VDD E net58 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD RB net13 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP11 net13 net79 net61 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net20 E net13 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP4 VDD CK net0301 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD net0301 net79 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net61 net90 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP13 net35 net90 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net35 net0301 net61 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net90 net0301 net37 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP16 VDD net37 net97 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD net97 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP29 net75 net97 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net75 net79 net37 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net53 D net13 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD net58 net53 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MN16 net58 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 net61 net0301 net73 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN11 net71 RB VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net73 net58 net77 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net70 E net71 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net73 D net70 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN17 net71 net75 net77 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 net0301 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net79 net0301 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net90 net61 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN12 net61 net79 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net90 net92 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net37 net79 net90 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN15 net97 net37 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN18 Q net97 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN25 net37 net0301 net75 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN29 VSS net97 net75 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
.ends DFEQZRM8HM
                                                           
.subckt DFERM1HM Q QB CK D E RB VDD VSS 
MN17 net46 net68 VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN6 net11 RB VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN16 net11 net13 net68 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN10 Q net68 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net46 net0193 net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 QB net46 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN13 net33 net62 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net0193 net44 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net35 net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net35 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net13 net62 net31 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net0182 E net44 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net44 net0185 net47 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net47 net46 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0182 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net0185 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net31 net29 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net62 net0193 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0193 CK VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP20 net31 net0193 net13 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 VDD RB net68 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP16 net68 net13 VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP15 VDD net68 net46 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP14 VDD net68 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP12 net13 net62 net46 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net46 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 net89 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net89 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net46 net96 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net96 E net99 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net99 net0185 net0182 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net29 net62 net99 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP7 VDD D net0182 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP8 VDD E net0185 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD net29 net31 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP11 net89 net0193 net29 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0193 net62 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP4 VDD CK net0193 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFERM1HM
                                                           
.subckt DFERM2HM Q QB CK D E RB VDD VSS 
MN17 net46 net68 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net11 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN16 net11 net13 net68 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN10 Q net68 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN15 net46 net0193 net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 QB net46 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN13 net33 net62 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net0193 net44 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN11 net35 net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net35 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net13 net62 net31 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net0182 E net44 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN3 net44 net0185 net47 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net47 net46 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net0182 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net0185 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net31 net29 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net62 net0193 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0193 CK VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP20 net31 net0193 net13 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 VDD RB net68 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP16 net68 net13 VDD VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 VDD net68 net46 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 VDD net68 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 net13 net62 net46 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net46 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 net89 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net89 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net46 net96 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP3 net96 E net99 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP5 net99 net0185 net0182 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net29 net62 net99 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP7 VDD D net0182 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD E net0185 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net29 net31 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP11 net89 net0193 net29 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0193 net62 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0193 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFERM2HM
                                                           
.subckt DFERM4HM Q QB CK D E RB VDD VSS 
MN17 net46 net68 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net11 RB VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN16 net11 net13 net68 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN10 Q net68 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN15 net46 net0193 net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 QB net46 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN13 net33 net62 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net0193 net44 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN11 net35 net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net35 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net13 net62 net31 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net0182 E net44 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN3 net44 net0185 net47 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net47 net46 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net0182 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net0185 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net31 net29 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net62 net0193 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0193 CK VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MP20 net31 net0193 net13 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 VDD RB net68 VDD P_15_LL_EE2_UCFN w=0.96u l=0.12u
MP16 net68 net13 VDD VDD P_15_LL_EE2_UCFN w=0.96u l=0.12u
MP15 VDD net68 net46 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 VDD net68 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP12 net13 net62 net46 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net46 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 net89 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net89 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net46 net96 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP3 net96 E net99 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP5 net99 net0185 net0182 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net29 net62 net99 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP7 VDD D net0182 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD E net0185 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net29 net31 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP11 net89 net0193 net29 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0193 net62 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0193 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFERM4HM
                                                           
.subckt DFERM8HM Q QB CK D E RB VDD VSS 
MN17 net46 net68 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN6 net11 RB VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN16 net11 net13 net68 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN10 Q net68 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN15 net46 net0193 net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 QB net46 VSS VSS N_15_LL_EE2_UCFN w=2.18u l=0.12u
MN13 net33 net62 net29 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net0193 net44 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN11 net35 net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net35 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net13 net62 net31 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net0182 E net44 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN3 net44 net0185 net47 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net47 net46 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net0182 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net0185 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net31 net29 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net62 net0193 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net0193 CK VSS VSS N_15_LL_EE2_UCFN w=0.4u l=0.12u
MP20 net31 net0193 net13 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP17 VDD RB net68 VDD P_15_LL_EE2_UCFN w=0.96u l=0.12u
MP16 net68 net13 VDD VDD P_15_LL_EE2_UCFN w=0.96u l=0.12u
MP15 VDD net68 net46 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP14 VDD net68 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP12 net13 net62 net46 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net46 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 net89 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 VDD RB net89 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net46 net96 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net96 E net99 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 net99 net0185 net0182 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net29 net62 net99 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP7 VDD D net0182 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP8 VDD E net0185 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net29 net31 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP11 net89 net0193 net29 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0193 net62 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP4 VDD CK net0193 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
.ends DFERM8HM
                                                           
.subckt DFEZRM1HM Q QB CK D E RB VDD VSS 
MP27 net0158 net11 net0135 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP24 net0118 D net0135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP23 VDD net0130 net0118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net0136 E net0135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD net079 net0136 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MN26 net0196 net079 net0184 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 VSS RB net0196 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN20 net0158 net050 net0192 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0192 D net0195 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN22 net0192 net0130 net0184 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN23 net0195 E net0196 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends DFEZRM1HM
                                                           
.subckt DFEZRM2HM Q QB CK D E RB VDD VSS 
MP27 net0158 net0227 net0135 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP24 net0118 D net0135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP23 VDD net0130 net0118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net0136 E net0135 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP21 VDD net079 net0136 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP14 net0128 net0227 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net0227 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MN26 net0196 net079 net0184 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN27 VSS RB net0196 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN20 net0158 net050 net0192 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0192 D net0195 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 net0192 net0130 net0184 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN23 net0195 E net0196 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 net019 net0227 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0227 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0227 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFEZRM2HM
                                                           
.subckt DFEZRM4HM Q QB CK D E RB VDD VSS 
MP27 net0158 net0228 net0135 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP24 net0118 D net0135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP23 VDD net0130 net0118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net0136 E net0135 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP21 VDD net079 net0136 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net0228 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.42u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.42u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net0228 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MN26 net0196 net079 net0184 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN27 VSS RB net0196 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN20 net0158 net050 net0192 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0192 D net0195 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 net0192 net0130 net0184 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN23 net0195 E net0196 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN8 net019 net0228 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0228 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0228 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFEZRM4HM
                                                           
.subckt DFEZRM8HM Q QB CK D E RB VDD VSS 
MP27 net0158 net0227 net0135 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP24 net0118 D net0135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP23 VDD net0130 net0118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net0136 E net0135 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP21 VDD net079 net0136 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.9u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=1.28u l=0.12u
MP14 net0128 net0227 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.44u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.48u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP16 VDD E net0130 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP8 VDD net0158 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net0158 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net0227 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MN26 net0196 net079 net0184 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN27 VSS RB net0196 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net0130 E VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN20 net0158 net050 net0192 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0192 D net0195 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 net0192 net0130 net0184 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN23 net0195 E net0196 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN8 net019 net0227 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net019 net0158 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net0158 net0227 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net0227 net050 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFEZRM8HM
                                                           
.subckt DFM1HM Q QB CK D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFM1HM
                                                           
.subckt DFM2HM Q QB CK D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFM2HM
                                                           
.subckt DFM4HM Q QB CK D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFM4HM
                                                           
.subckt DFM8HM Q QB CK D VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFM8HM
                                                           
.subckt DFMM1HM Q QB CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN30 QB net48 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP30 VDD net48 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFMM1HM
                                                           
.subckt DFMM2HM Q QB CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN30 QB net48 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP30 VDD net48 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFMM2HM
                                                           
.subckt DFMM4HM Q QB CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN30 QB net48 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=1.26u l=0.12u
MP30 VDD net48 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=1.26u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFMM4HM
                                                           
.subckt DFMM8HM Q QB CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN30 QB net48 VSS VSS N_15_LL_EE2_UCFN w=2.18u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=1.48u l=0.12u
MP30 VDD net48 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=2.96u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=1.24u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
.ends DFMM8HM
                                                           
.subckt DFMQM1HM Q CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFMQM1HM
                                                           
.subckt DFMQM2HM Q CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFMQM2HM
                                                           
.subckt DFMQM4HM Q CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=1.26u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=1.26u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
.ends DFMQM4HM
                                                           
.subckt DFMQM8HM Q CK D1 D2 S VDD VSS 
MN9 net0130 S VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0133 D2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net20 net0285 net15 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 net17 D1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net20 S net17 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0133 net0130 net20 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN10 net31 net15 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN12 net15 net56 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 VSS net31 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net86 net56 net31 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net38 net86 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN18 Q net38 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN25 net86 net0285 net48 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 VSS net38 net48 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net56 net0285 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN4 net0285 CK VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP8 VDD S net0130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D2 net0133 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP6 net15 net56 net69 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net69 S net0133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net72 net0130 net69 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD D1 net72 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net15 net31 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP13 net84 net31 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net84 net0285 net15 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net31 net0285 net86 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 VDD net86 net38 VDD P_15_LL_EE2_UCFN w=1.48u l=0.12u
MP19 VDD net38 Q VDD P_15_LL_EE2_UCFN w=2.96u l=0.12u
MP29 net48 net38 VDD VDD P_15_LL_EE2_UCFN w=1.24u l=0.12u
MP26 net48 net56 net86 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net0285 net56 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP4 VDD CK net0285 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
.ends DFMQM8HM
                                                           
.subckt DFQM1HM Q CK D VDD VSS 
MP16 net078 net050 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 net078 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP9 net0128 net11 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net11 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net11 net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net050 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN16 net0128 net11 net0114 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net019 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN15 VSS net0124 net0114 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net050 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net11 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net050 net11 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net11 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFQM1HM
                                                           
.subckt DFQM2HM Q CK D VDD VSS 
MP16 net085 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 net085 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN16 net0128 net050 net080 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 VSS net0124 net080 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQM2HM
                                                           
.subckt DFQM4HM Q CK D VDD VSS 
MP16 net088 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 net088 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN15 VSS net0124 net080 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net0128 net050 net080 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQM4HM
                                                           
.subckt DFQM8HM Q CK D VDD VSS 
MP16 net085 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 net085 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN15 VSS net0124 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net0128 net050 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFQM8HM
                                                           
.subckt DFQRM1HM Q CK D RB VDD VSS 
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0102 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0102 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net0128 net050 net090 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 VSS net0124 net090 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQRM1HM
                                                           
.subckt DFQRM2HM Q CK D RB VDD VSS 
MP18 net0145 RB VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP24 net0102 net0145 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0102 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0145 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0145 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net0128 net050 net089 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 VSS net0145 net089 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0145 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN15 net0145 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQRM2HM
                                                           
.subckt DFQRM4HM Q CK D RB VDD VSS 
MP18 net0145 RB VDD VDD P_15_LL_EE2_UCFN w=0.8u l=0.12u
MP24 net0102 net0145 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0102 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0145 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0145 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net0128 net050 net089 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 VSS net0145 net089 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0145 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN15 net0145 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQRM4HM
                                                           
.subckt DFQRM8HM Q CK D RB VDD VSS 
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.8u l=0.12u
MP24 net0102 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0102 net11 net0128 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.06u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net0128 net050 net090 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 VSS net0124 net090 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
.ends DFQRM8HM
                                                           
.subckt DFQRSM1HM Q CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQRSM1HM
                                                           
.subckt DFQRSM2HM Q CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQRSM2HM
                                                           
.subckt DFQRSM4HM Q CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFQRSM4HM
                                                           
.subckt DFQRSM8HM Q CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=1u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
.ends DFQRSM8HM
                                                           
.subckt DFQSM1HM Q CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends DFQSM1HM
                                                           
.subckt DFQSM2HM Q CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFQSM2HM
                                                           
.subckt DFQSM4HM Q CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFQSM4HM
                                                           
.subckt DFQSM8HM Q CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
.ends DFQSM8HM
                                                           
.subckt DFQZRM1HM Q CK D RB VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFQZRM1HM
                                                           
.subckt DFQZRM2HM Q CK D RB VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFQZRM2HM
                                                           
.subckt DFQZRM4HM Q CK D RB VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFQZRM4HM
                                                           
.subckt DFQZRM8HM Q CK D RB VDD VSS 
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFQZRM8HM
                                                           
.subckt DFRM1HM Q QB CK D RB VDD VSS 
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFRM1HM
                                                           
.subckt DFRM2HM Q QB CK D RB VDD VSS 
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFRM2HM
                                                           
.subckt DFRM4HM Q QB CK D RB VDD VSS 
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.79u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.90u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFRM4HM
                                                           
.subckt DFRM8HM Q QB CK D RB VDD VSS 
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.79u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.86u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2.18u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
.ends DFRM8HM
                                                           
.subckt DFRSM1HM Q QB CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends DFRSM1HM
                                                           
.subckt DFRSM2HM Q QB CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFRSM2HM
                                                           
.subckt DFRSM4HM Q QB CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.85u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.01u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFRSM4HM
                                                           
.subckt DFRSM8HM Q QB CK D RB SB VDD VSS 
MP20 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net0124 RB VDD VDD P_15_LL_EE2_UCFN w=0.85u l=0.12u
MP23 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP22 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP19 VDD RB net024 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.01u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN24 net0164 SB net019 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN23 net0164 net047 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN18 VSS RB net0142 VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2.18u l=0.12u
MN21 net079 SB net0171 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN17 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN22 VSS net0124 net0171 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net0124 net0128 net0142 VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN6 net0147 net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
.ends DFRSM8HM
                                                           
.subckt DFSM1HM Q QB CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFSM1HM
                                                           
.subckt DFSM2HM Q QB CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFSM2HM
                                                           
.subckt DFSM4HM Q QB CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.6u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFSM4HM
                                                           
.subckt DFSM8HM Q QB CK D SB VDD VSS 
MP20 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SB net079 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP16 net019 SB VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.2u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP5 net027 D net047 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD net11 net027 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN18 net079 SB net0144 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN17 VSS net0124 net0144 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN15 net0152 SB net019 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN16 net0152 net047 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.6u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net044 net050 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN3 net047 D net044 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
.ends DFSM8HM
                                                           
.subckt DFZRM1HM Q QB CK D RB VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFZRM1HM
                                                           
.subckt DFZRM2HM Q QB CK D RB VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFZRM2HM
                                                           
.subckt DFZRM4HM Q QB CK D RB VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.32u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends DFZRM4HM
                                                           
.subckt DFZRM8HM Q QB CK D RB VDD VSS 
MP15 VDD net079 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 net079 net0124 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP14 net0128 net11 net079 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD net0124 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net0128 net0124 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0128 net050 net019 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 VDD net047 net019 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP7 net024 net050 net047 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 net024 net019 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 VDD net050 net11 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net027 net11 net047 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD D net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD CK net050 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP16 VDD RB net027 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MN14 QB net079 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN12 VSS net0124 net079 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net079 net050 net0128 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 Q net0124 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN9 net0124 net0128 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN8 net019 net11 net0128 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net019 net047 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 VSS net019 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net047 net11 net039 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net0136 RB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net044 D net0136 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net11 net050 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net047 net050 net044 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net050 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends DFZRM8HM
                                                           
.subckt FIL16HM VDD VSS
.ends FIL16HM
                                                           
.subckt FIL1HM VDD VSS
.ends FIL1HM
                                                           
.subckt FIL2HM VDD VSS
.ends FIL2HM
                                                           
.subckt FIL32HM VDD VSS
.ends FIL32HM
                                                           
.subckt FIL4HM VDD VSS
.ends FIL4HM
                                                           
.subckt FIL64HM VDD VSS
.ends FIL64HM
                                                           
.subckt FIL8HM VDD VSS
.ends FIL8HM
                                                           
.subckt FILE128HM VDD VSS 
MN0 VSS net02 net02 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 VSS net04 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=2.70u
MP0 VDD net01 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net04 net02 VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 VDD net03 VDD VDD P_15_LL_EE2_UCFN w=7.68u l=2.70u
.ends FILE128HM
                                                           
.subckt FILE16HM VDD VSS 
MN0 VSS net02 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 VSS net04 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=2.04u
MP0 VDD net01 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net04 net02 VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 VDD net03 VDD VDD P_15_LL_EE2_UCFN w=0.96u l=2.04u
.ends FILE16HM
                                                           
.subckt FILE32HM VDD VSS 
MN0 VSS net02 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN2 VSS net04 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=2.42u
MP0 VDD net01 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net04 net02 VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 VDD net03 VDD VDD P_15_LL_EE2_UCFN w=1.92u l=2.42u
.ends FILE32HM
                                                           
.subckt FILE3HM VDD VSS 
MN0 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.32u
MP0 net01 net02 VDD VDD P_15_LL_EE2_UCFN w=0.54u l=0.32u
.ends FILE3HM
                                                           
.subckt FILE4HM VDD VSS 
MN0 VSS net01 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.20u
MN1 VSS net01 net02 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MP0 VDD net02 VDD VDD P_15_LL_EE2_UCFN w=0.54u l=0.20u
MP1 VDD net02 net01 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
.ends FILE4HM
                                                           
.subckt FILE64HM VDD VSS 
MN0 VSS net02 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN2 VSS net04 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=2.61u
MP0 VDD net01 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net04 net02 VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 VDD net03 VDD VDD P_15_LL_EE2_UCFN w=3.84u l=2.61u
.ends FILE64HM
                                                           
.subckt FILE8HM VDD VSS 
MN0 VSS net02 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN2 VSS net04 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=1.28u
MP0 VDD net01 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net04 net02 VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 VDD net03 VDD VDD P_15_LL_EE2_UCFN w=0.48u l=1.28u
.ends FILE8HM
                                                           
.subckt INVM0HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends INVM0HM
                                                           
.subckt INVM10HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.80u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=3.40u l=0.12u
.ends INVM10HM
                                                           
.subckt INVM12HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends INVM12HM
                                                           
.subckt INVM14HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=3.92u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=4.76u l=0.12u
.ends INVM14HM
                                                           
.subckt INVM16HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends INVM16HM
                                                           
.subckt INVM18HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=5.04u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=6.12u l=0.12u
.ends INVM18HM
                                                           
.subckt INVM1HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends INVM1HM
                                                           
.subckt INVM20HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=5.60u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=6.80u l=0.12u
.ends INVM20HM
                                                           
.subckt INVM24HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=6.72u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
.ends INVM24HM
                                                           
.subckt INVM28HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=7.84u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=9.52u l=0.12u
.ends INVM28HM
                                                           
.subckt INVM2HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends INVM2HM
                                                           
.subckt INVM32HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=8.96u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
.ends INVM32HM
                                                           
.subckt INVM36HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=10.08u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=12.24u l=0.12u
.ends INVM36HM
                                                           
.subckt INVM3HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
.ends INVM3HM
                                                           
.subckt INVM40HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=10.64u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=12.92u l=0.12u
.ends INVM40HM
                                                           
.subckt INVM48HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=12.88u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=15.64u l=0.12u
.ends INVM48HM
                                                           
.subckt INVM4HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends INVM4HM
                                                           
.subckt INVM5HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.41u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.71u l=0.12u
.ends INVM5HM
                                                           
.subckt INVM6HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends INVM6HM
                                                           
.subckt INVM8HM Z A VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends INVM8HM
                                                           
.subckt LACM0HM Q QB D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACM0HM
                                                           
.subckt LACM1HM Q QB D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACM1HM
                                                           
.subckt LACM2HM Q QB D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACM2HM
                                                           
.subckt LACM4HM Q QB D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACM4HM
                                                           
.subckt LACQM0HM Q D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACQM0HM
                                                           
.subckt LACQM1HM Q D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACQM1HM
                                                           
.subckt LACQM2HM Q D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACQM2HM
                                                           
.subckt LACQM4HM Q D GB VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 GB VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net12 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN0 net45 net15 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD GB net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net52 net12 net45 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net55 net15 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LACQM4HM
                                                           
.subckt LACQRSM0HM Q D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LACQRSM0HM
                                                           
.subckt LACQRSM1HM Q D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LACQRSM1HM
                                                           
.subckt LACQRSM2HM Q D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends LACQRSM2HM
                                                           
.subckt LACQRSM4HM Q D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends LACQRSM4HM
                                                           
.subckt LACRSM0HM Q QB D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LACRSM0HM
                                                           
.subckt LACRSM1HM Q QB D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LACRSM1HM
                                                           
.subckt LACRSM2HM Q QB D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends LACRSM2HM
                                                           
.subckt LACRSM4HM Q QB D GB RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN8 net19 GB VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 GB net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 net19 net49 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD GB net19 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 net19 net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net65 GB net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends LACRSM4HM
                                                           
.subckt LAGCEM12HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=1.5u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=1.46u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=1.77u l=0.12u
.ends LAGCEM12HM
                                                           
.subckt LAGCEM16HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=1.41u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=1.41u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=1.90u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=2.36u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=2.32u l=0.12u
.ends LAGCEM16HM
                                                           
.subckt LAGCEM20HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=1.76u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=1.76u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=2.5u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=2.54u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.66u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=2.37u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=6.80u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=6.80u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=2.36u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=3.40u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.81u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=2.90u l=0.12u
.ends LAGCEM20HM
                                                           
.subckt LAGCEM2HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
.ends LAGCEM2HM
                                                           
.subckt LAGCEM3HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
.ends LAGCEM3HM
                                                           
.subckt LAGCEM4HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
.ends LAGCEM4HM
                                                           
.subckt LAGCEM6HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=0.76u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=1.96u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=1.96u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=0.90u l=0.12u
.ends LAGCEM6HM
                                                           
.subckt LAGCEM8HM GCK CK E VDD VSS 
MN8 GCK net2 VSS VSS N_15_LL_EE2_UCFN w=0.69u l=0.12u
MN7 GCK net16 VSS VSS N_15_LL_EE2_UCFN w=0.69u l=0.12u
MN6 net076 net2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net14 E VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN4 net2 net16 net14 VSS N_15_LL_EE2_UCFN w=0.98u l=0.12u
MN3 VSS net076 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net2 net5 net12 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net5 net16 VSS VSS N_15_LL_EE2_UCFN w=0.30u l=0.12u
MN0 net16 CK VSS VSS N_15_LL_EE2_UCFN w=1.00u l=0.12u
MP7 VDD net16 net072 VDD P_15_LL_EE2_UCFN w=2.64u l=0.12u
MP8 net072 net2 GCK VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP6 VDD net2 net076 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP5 net36 net076 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 net36 net16 net2 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 net39 net5 net2 VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
MP2 VDD E net39 VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP1 VDD net16 net5 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD CK net16 VDD P_15_LL_EE2_UCFN w=1.22u l=0.12u
.ends LAGCEM8HM

.subckt LAGCECSM12HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=1.35u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=1.35u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=1.7u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends LAGCECSM12HM
                                                           
.subckt LAGCECSM16HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=1.8u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=1.8u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=2.225u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends LAGCECSM16HM
                                                           
.subckt LAGCECSM20HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=2.25u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=2.25u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=2.91u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=3.4u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=3.4u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=6.8u l=0.12u
.ends LAGCECSM20HM
                                                           
.subckt LAGCECSM2HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends LAGCECSM2HM
                                                           
.subckt LAGCECSM3HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
.ends LAGCECSM3HM
                                                           
.subckt LAGCECSM4HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends LAGCECSM4HM
                                                           
.subckt LAGCECSM6HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=0.68u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=0.68u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.86u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends LAGCECSM6HM
                                                           
.subckt LAGCECSM8HM GCK CKB E SE VDD VSS 
MN11 net0178 net32 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN10 net30 CKB VSS VSS N_15_LL_EE2_UCFN w=0.90u l=0.12u
MN9 net30 net0178 VSS VSS N_15_LL_EE2_UCFN w=0.90u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net57 CKB VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net54 net57 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=1.14u l=0.12u
MP11 VDD net32 net0178 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net0178 net0179 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 net0179 CKB net30 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CKB net57 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net57 net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends LAGCECSM8HM
                                                          
.subckt LAGCESM12HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.64u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.64u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=1.7u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends LAGCESM12HM
                                                           
.subckt LAGCESM16HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.86u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.86u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=2.28u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=5.48u l=0.12u
.ends LAGCESM16HM
                                                           
.subckt LAGCESM20HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=2.88u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=1.71u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=1.71u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=6.84u l=0.12u
.ends LAGCESM20HM
                                                           
.subckt LAGCESM2HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends LAGCESM2HM
                                                           
.subckt LAGCESM3HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
.ends LAGCESM3HM
                                                           
.subckt LAGCESM4HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends LAGCESM4HM
                                                           
.subckt LAGCESM6HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=0.86u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends LAGCESM6HM
                                                           
.subckt LAGCESM8HM GCK CK E SE VDD VSS 
MN10 net6 CK VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN9 net30 net32 net6 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 net32 net24 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net54 CK VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN6 net57 net54 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 VSS net32 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net24 net57 net16 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net21 SE VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net21 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net24 net54 net21 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 GCK net30 VSS VSS N_15_LL_EE2_UCFN w=1.14u l=0.12u
MP10 VDD net32 net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 VDD CK net30 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD net24 net32 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD CK net54 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP6 VDD net54 net57 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net37 net32 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 net37 net54 net24 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net40 E net46 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SE net40 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net46 net57 net24 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net30 GCK VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends LAGCESM8HM
                                                           
.subckt LAM0HM Q QB D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAM0HM
                                                           
.subckt LAM1HM Q QB D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAM1HM
                                                           
.subckt LAM2HM Q QB D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAM2HM
                                                           
.subckt LAM4HM Q QB D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 QB net56 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD net56 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAM4HM
                                                           
.subckt LAQM0HM Q D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAQM0HM
                                                           
.subckt LAQM1HM Q D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAQM1HM
                                                           
.subckt LAQM2HM Q D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAQM2HM
                                                           
.subckt LAQM4HM Q D G VDD VSS 
MN8 Q net45 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net56 net45 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net12 net15 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net15 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net36 net56 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net45 net15 net36 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net42 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net45 net12 net42 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 VDD net45 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP7 VDD net45 net56 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net15 net12 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD G net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D net52 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net52 net15 net45 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net55 net12 net45 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net56 net55 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends LAQM4HM
                                                           
.subckt LAQRSM0HM Q D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LAQRSM0HM
                                                           
.subckt LAQRSM1HM Q D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LAQRSM1HM
                                                           
.subckt LAQRSM2HM Q D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends LAQRSM2HM
                                                           
.subckt LAQRSM4HM Q D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends LAQRSM4HM
                                                           
.subckt LARSM0HM Q QB D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LARSM0HM
                                                           
.subckt LARSM1HM Q QB D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends LARSM1HM
                                                           
.subckt LARSM2HM Q QB D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends LARSM2HM
                                                           
.subckt LARSM4HM Q QB D G RB SB VDD VSS 
MN9 net094 net64 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net13 net54 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN10 QB net54 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN7 net54 SB net094 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN8 net19 G VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 Q net13 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN5 net37 net54 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net37 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net64 net19 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN1 net49 D net46 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN0 net64 G net49 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MP10 VDD net54 net13 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP6 VDD net64 net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP9 VDD net54 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP8 VDD SB net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP7 VDD G net19 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD net13 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net59 net54 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP3 net59 G net64 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 net65 net19 net64 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD D net65 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends LARSM4HM
                                                           
.subckt MAO222M0HM Z A B C VDD VSS 
MN0 net03 A VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN1 net01 A net05 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN2 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN4 net01 C net03 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP1 net04 A net01 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net02 C net01 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends MAO222M0HM
                                                           
.subckt MAO222M1HM Z A B C VDD VSS 
MN0 net03 A VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN1 net01 A net05 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN2 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN4 net01 C net03 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP1 net04 A net01 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net02 C net01 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends MAO222M1HM
                                                           
.subckt MAO222M2HM Z A B C VDD VSS 
MN0 net03 A VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN1 net01 A net05 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN2 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN3 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN4 net01 C net03 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP1 net04 A net01 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net02 C net01 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MAO222M2HM
                                                           
.subckt MAO222M4HM Z A B C VDD VSS 
MN0 net01 A net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net01 A net03 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN5 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net04 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net05 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net04 B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MAO222M4HM
                                                           
.subckt MAOI2223M0HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN3 Z D net01 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN4 Z A net02 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN5 net02 B net03 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN6 net03 C VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP3 net04 D Z VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP4 net05 A Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 net06 B net05 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP6 VDD C net06 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends MAOI2223M0HM
                                                           
.subckt MAOI2223M1HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z D net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z A net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN5 net02 B net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN6 net03 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP3 net04 D Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP4 net05 A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 net06 B net05 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP6 VDD C net06 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends MAOI2223M1HM
                                                           
.subckt MAOI2223M2HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 Z D net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 Z A net02 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN5 net02 B net03 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN6 net03 C VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MP0 VDD A net04 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP1 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP2 VDD C net04 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP3 net04 D Z VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP4 net05 A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net06 B net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD C net06 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MAOI2223M2HM
                                                           
.subckt MAOI2223M4HM Z A B C D VDD VSS 
MN0 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net01 D net02 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net01 A net03 VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN5 net03 B net04 VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN6 net04 C VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN7 net08 net01 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN8 Z net08 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net05 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP1 VDD B net05 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP2 VDD C net05 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP3 net05 D net01 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP4 net06 A net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net07 B net06 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP6 VDD C net07 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD net01 net08 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 VDD net08 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MAOI2223M4HM
                                                           
.subckt MAOI222M0HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN1 Z A net02 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN2 Z B net01 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN3 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MP0 net03 A Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net04 A Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net03 B Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends MAOI222M0HM
                                                           
.subckt MAOI222M1HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 Z A net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 Z B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 net03 A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net04 A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net03 B Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends MAOI222M1HM
                                                           
.subckt MAOI222M2HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN1 Z A net02 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN2 Z B net01 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN3 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 net03 A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net04 A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MAOI222M2HM
                                                           
.subckt MAOI222M4HM Z A B C VDD VSS 
MN0 net05 A net01 VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN1 net05 A net02 VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN2 net05 B net01 VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN3 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN5 net06 net05 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN6 Z net06 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A net05 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net04 A net05 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 net03 B net05 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD B net04 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 VDD net05 net06 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 VDD net06 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MAOI222M4HM
                                                           
.subckt MAOI22M0HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MP0 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP1 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP2 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net04 A2 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends MAOI22M0HM
                                                           
.subckt MAOI22M1HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MP0 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP1 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP2 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net04 A2 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends MAOI22M1HM
                                                           
.subckt MAOI22M2HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN3 net03 A2 VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.4u l=0.12u
MP0 net02 B1 net01 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP1 VDD B2 net02 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP2 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net04 A2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MAOI22M2HM
                                                           
.subckt MAOI22M4HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 net02 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net03 B1 net04 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN3 net03 B2 net04 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN4 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A1 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD A2 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MAOI22M4HM
                                                           
.subckt MOAI22M0HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 B1 net02 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 Z A2 net03 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
.ends MOAI22M0HM
                                                           
.subckt MOAI22M1HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 B1 net02 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 Z A2 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.30u l=0.12u
.ends MOAI22M1HM
                                                           
.subckt MOAI22M2HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 B1 net02 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN3 Z A2 net03 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN4 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD B1 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD B2 net01 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends MOAI22M2HM
                                                           
.subckt MOAI22M4HM Z A1 A2 B1 B2 VDD VSS 
MN0 net01 A1 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net03 B1 net04 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN3 net04 B2 VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN4 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A1 net01 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net05 B2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MOAI22M4HM
                                                           
.subckt MUX2M0HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
.ends MUX2M0HM
                                                           
.subckt MUX2M1HM Z A B S VDD VSS 
MN5 net30 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net04 net30 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net02 S net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 net30 S VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 net11 A VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 net11 S net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 net12 net30 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net12 B VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 Z net01 VDD VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends MUX2M1HM
                                                           
.subckt MUX2M2HM Z A B S VDD VSS 
MN5 net30 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net04 net30 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net02 S net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP5 net30 S VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP4 net11 A VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 net11 S net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 net12 net30 net01 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net12 B VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 Z net01 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MUX2M2HM
                                                           
.subckt MUX2M3HM Z A B S VDD VSS 
MN5 net30 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 A VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net04 net30 net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 S net01 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN0 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MP5 net30 S VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP4 net11 A VDD VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP3 net11 S net01 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP2 net12 net30 net01 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 net12 B VDD VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 Z net01 VDD VDD P_15_LL_EE2_UCFN w=1.02u l=0.12u
.ends MUX2M3HM
                                                           
.subckt MUX2M4HM Z A B S VDD VSS 
MN5 net30 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 A VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN3 net04 net30 net01 VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN2 net02 S net01 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.50u l=0.12u
MN0 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP5 net30 S VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP4 net11 A VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP3 net11 S net01 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 net12 net30 net01 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP1 net12 B VDD VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 Z net01 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MUX2M4HM
                                                           
.subckt MUX2M6HM Z A B S VDD VSS 
MN5 net30 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 A VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN3 net04 net30 net01 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN2 net02 S net01 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP5 net30 S VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP4 net11 A VDD VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP3 net11 S net01 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 net12 net30 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net12 B VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 Z net01 VDD VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends MUX2M6HM
                                                           
.subckt MUX2M8HM Z A B S VDD VSS 
MN5 Z net10 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN4 net18 S net10 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net15 S VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net18 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP5 VDD net10 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 net10 net15 net18 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP2 VDD S net15 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net10 S net071 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP1 VDD B net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MUX2M8HM
                                                           
.subckt MUX3M0HM Z A B C S0 S1 VDD VSS 
MN9 net01 S0 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net02 net01 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN6 net03 S0 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN5 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net04 S1 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net05 net04 net11 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net06 S1 net11 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net06 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net11 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP9 net01 S0 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net07 A VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP7 net07 S0 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP6 net08 net01 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP5 net08 B VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP4 net04 S1 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 net09 S1 net11 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 net10 net04 net11 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 net10 C VDD VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP0 Z net11 VDD VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends MUX3M0HM
                                                           
.subckt MUX3M1HM Z A B C S0 S1 VDD VSS 
MN9 net01 S0 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net02 net01 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN6 net03 S0 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN5 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net04 S1 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net05 net04 net11 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net06 S1 net11 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net06 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net11 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 net01 S0 VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP8 net07 A VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP7 net07 S0 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP6 net08 net01 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP5 net08 B VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP4 net04 S1 VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP3 net09 S1 net11 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 net10 net04 net11 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 net10 C VDD VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP0 Z net11 VDD VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends MUX3M1HM
                                                           
.subckt MUX3M2HM Z A B C S0 S1 VDD VSS 
MN9 net01 S0 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net02 net01 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN6 net03 S0 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN5 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net04 S1 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net05 net04 net11 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net06 S1 net11 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net06 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net11 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP9 net01 S0 VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP8 net07 A VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP7 net07 S0 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP6 net08 net01 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP5 net08 B VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP4 net04 S1 VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP3 net09 S1 net11 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 net10 net04 net11 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP1 net10 C VDD VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP0 Z net11 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MUX3M2HM
                                                           
.subckt MUX3M4HM Z A B C S0 S1 VDD VSS 
MN9 net01 S0 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN7 net02 net01 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN6 net03 S0 net05 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN5 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net04 S1 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net05 net04 net11 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN2 net06 S1 net11 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN1 net06 C VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN0 Z net11 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP9 net01 S0 VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP8 net07 A VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP7 net07 S0 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP6 net08 net01 net09 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP5 net08 B VDD VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP4 net04 S1 VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP3 net09 S1 net11 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP2 net10 net04 net11 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 net10 C VDD VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 Z net11 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends MUX3M4HM
                                                           
.subckt MUX4M0HM Z A B C D S0 S1 VDD VSS 
MN18 net098 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net082 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net098 S0 net0108 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN22 net0110 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net15 S0 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net065 S1 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0110 net15 net0108 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN26 net10 S1 net0120 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net082 S0 net10 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net0108 net065 net0120 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 Z net0120 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net071 C VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP27 net0120 S1 net0108 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net10 net15 net082 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 net0108 net15 net098 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD S1 net065 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD B net098 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net0108 S0 net0110 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 VDD A net0110 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD S0 net15 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP26 net0120 net065 net10 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D net082 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net10 S0 net071 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD net0120 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP0 VDD C net071 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends MUX4M0HM
                                                           
.subckt MUX4M1HM Z A B C D S0 S1 VDD VSS 
MN18 net098 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net082 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net098 S0 net0108 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN22 net0110 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net15 S0 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net065 S1 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0110 net15 net0108 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN26 net10 S1 net0120 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net082 S0 net10 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net0108 net065 net0120 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 Z net0120 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN0 net071 C VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP27 net0120 S1 net0108 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net10 net15 net082 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 net0108 net15 net098 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD S1 net065 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD B net098 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net0108 S0 net0110 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 VDD A net0110 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD S0 net15 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP26 net0120 net065 net10 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD D net082 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net10 S0 net071 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD net0120 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP0 VDD C net071 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends MUX4M1HM
                                                           
.subckt MUX4M2HM Z A B C D S0 S1 VDD VSS 
MN18 net098 B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN7 net082 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN21 net098 S0 net0108 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN22 net0110 A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN10 net15 S0 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN19 net065 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN20 net0110 net15 net0108 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN26 net10 S1 net0120 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net082 S0 net10 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN27 net0108 net065 net0120 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN17 Z net0120 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net071 C VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP27 net0120 S1 net0108 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net10 net15 net082 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP18 net0108 net15 net098 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD S1 net065 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP20 VDD B net098 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP21 net0108 S0 net0110 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP22 VDD A net0110 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP10 VDD S0 net15 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP26 net0120 net065 net10 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP7 VDD D net082 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 net10 S0 net071 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 VDD net0120 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD C net071 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
.ends MUX4M2HM
                                                           
.subckt MUX4M4HM Z A B C D S0 S1 VDD VSS 
MN18 net098 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net082 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net098 S0 net0108 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN22 net0110 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN10 net15 S0 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN19 net065 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN20 net0110 net15 net0108 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN26 net10 S1 net0120 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN3 net071 net15 net10 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN6 net082 S0 net10 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN27 net0108 net065 net0120 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN17 Z net0120 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN0 net071 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP27 net0120 S1 net0108 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP6 net10 net15 net082 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP18 net0108 net15 net098 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP19 VDD S1 net065 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP20 VDD B net098 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 net0108 S0 net0110 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP22 VDD A net0110 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD S0 net15 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP26 net0120 net065 net10 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP7 VDD D net082 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net10 S0 net071 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP17 VDD net0120 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP0 VDD C net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends MUX4M4HM
                                                           
.subckt MXB2M0HM Z A B S VDD VSS 
MP12 VDD B net70 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP13 net70 net75 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP11 VDD S net75 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 net64 S Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP14 VDD A net64 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MN11 net75 S VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN13 net84 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN14 Z S net78 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN15 net78 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN12 Z net75 net84 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends MXB2M0HM
                                                           
.subckt MXB2M1HM Z A B S VDD VSS 
MP12 VDD B net70 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP13 net70 net75 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP11 VDD S net75 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 net64 S Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP14 VDD A net64 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MN11 net75 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net84 A VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN14 Z S net78 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN15 net78 B VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN12 Z net75 net84 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends MXB2M1HM
                                                           
.subckt MXB2M2HM Z A B S VDD VSS 
MP12 VDD B net70 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net70 net75 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD S net75 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 net64 S Z VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP14 VDD A net64 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MN11 net75 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN13 net84 A VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN14 Z S net78 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN15 net78 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 Z net75 net84 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
.ends MXB2M2HM
                                                           
.subckt MXB2M3HM Z A B S VDD VSS 
MP6 VDD S net059 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP7 VDD A net056 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net21 Z VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP10 VDD net069 net21 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD B net062 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 net069 net059 net062 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 net069 S net056 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MN10 net21 net069 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net21 VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN7 net056 A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net059 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net062 B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net062 S net069 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net056 net059 net069 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends MXB2M3HM
                                                           
.subckt MXB2M4HM Z A B S VDD VSS 
MP6 VDD S net059 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP7 VDD A net056 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net21 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP10 VDD net069 net21 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD B net062 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP8 net069 net059 net062 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 net069 S net056 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MN10 net21 net069 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net056 A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net059 S VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net062 B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net062 S net069 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net056 net059 net069 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends MXB2M4HM
                                                           
.subckt MXB2M6HM Z A B S VDD VSS 
MP6 VDD S net059 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP7 VDD A net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net21 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP10 VDD net069 net21 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP5 VDD B net062 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP8 net069 net059 net062 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP9 net069 S net056 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MN10 net21 net069 VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN4 Z net21 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN7 net056 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net059 S VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net062 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net062 S net069 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN9 net056 net059 net069 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
.ends MXB2M6HM
                                                           
.subckt MXB2M8HM Z A B S VDD VSS 
MP6 VDD S net059 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP7 VDD A net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net21 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP10 VDD net069 net21 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD B net062 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP8 net069 net059 net062 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP9 net069 S net056 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MN10 net21 net069 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net21 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN7 net056 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net059 S VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net062 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net062 S net069 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN9 net056 net059 net069 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
.ends MXB2M8HM
                                                           
.subckt MXB3M0HM Z A B C S0 S1 VDD VSS 
MP14 net060 S0 net071 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net060 net068 net065 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD B net065 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP11 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP10 VDD S0 net068 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP6 VDD S1 net0127 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP7 VDD C net077 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP8 Z S1 net060 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP9 Z net0127 net077 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 net071 net068 net060 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN13 net065 S0 net060 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net065 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN11 net068 S0 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN10 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN7 net077 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN6 net0127 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net060 net0127 Z VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net077 S1 Z VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends MXB3M0HM
                                                           
.subckt MXB3M1HM Z A B C S0 S1 VDD VSS 
MP14 net060 S0 net071 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP13 net060 net068 net065 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD B net065 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD S0 net068 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP6 VDD S1 net0127 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP7 VDD C net077 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 Z S1 net060 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP9 Z net0127 net077 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MN14 net071 net068 net060 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN13 net065 S0 net060 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net065 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net068 S0 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN10 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net077 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net0127 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net060 net0127 Z VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net077 S1 Z VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends MXB3M1HM
                                                           
.subckt MXB3M2HM Z A B C S0 S1 VDD VSS 
MP14 net060 S0 net071 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP13 net060 net068 net065 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD B net065 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP10 VDD S0 net068 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP15 VDD net0190 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD S1 net0149 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP7 VDD C net077 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net087 net0190 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 net087 S1 net060 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP9 net087 net0149 net077 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MN15 Z net0190 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 net071 net068 net060 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN13 net065 S0 net060 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN12 net065 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net068 S0 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN10 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net0190 net087 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN7 net077 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN6 net0149 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net060 net0149 net087 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net077 S1 net087 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends MXB3M2HM
                                                           
.subckt MXB3M4HM Z A B C S0 S1 VDD VSS 
MP14 net060 S0 net071 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP13 net060 net068 net065 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD B net065 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP11 VDD A net071 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP10 VDD S0 net068 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP15 VDD net0190 Z VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MP6 VDD S1 net0149 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD C net077 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP4 VDD net087 net0190 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP8 net087 S1 net060 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP9 net087 net0149 net077 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MN15 Z net0190 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN14 net071 net068 net060 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN13 net065 S0 net060 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN12 net065 B VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN11 net068 S0 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN10 net071 A VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 net0190 net087 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN7 net077 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN6 net0149 S1 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 net060 net0149 net087 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN9 net077 S1 net087 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
.ends MXB3M4HM
                                                           
.subckt MXB4M0HM Z A B C D S0 S1 VDD VSS 
MP31 net177 S0 net178 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net184 S0 net198 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD A net177 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP23 net184 net201 net183 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP30 net180 net201 net178 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP26 VDD S1 net203 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP27 Z net203 net184 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 Z S1 net178 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD D net183 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP18 VDD C net198 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP20 VDD B net180 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP17 VDD S0 net201 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MN31 net178 net201 net177 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net198 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 net198 net201 net184 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN23 net183 S0 net184 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net177 A VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN30 net178 S0 net180 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN26 net203 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN27 net184 S1 Z VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net178 net203 Z VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net180 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN19 net183 D VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN17 net201 S0 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends MXB4M0HM
                                                           
.subckt MXB4M1HM Z A B C D S0 S1 VDD VSS 
MP29 net180 net201 net178 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP30 net177 S0 net178 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP22 net184 S0 net198 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP21 VDD A net177 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net184 net201 net183 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 VDD S1 net203 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP27 Z net203 net184 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP28 Z S1 net178 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD D net183 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP18 VDD C net198 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 VDD B net180 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP17 VDD S0 net201 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MN29 net178 S0 net180 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN18 net198 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 net198 net201 net184 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN23 net183 S0 net184 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN21 net177 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN30 net178 net201 net177 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN26 net203 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN27 net184 S1 Z VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN28 net178 net203 Z VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN20 net180 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 net183 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN17 net201 S0 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends MXB4M1HM
                                                           
.subckt MXB4M2HM Z A B C D S0 S1 VDD VSS 
MP32 net180 net201 net178 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP30 VDD net184 net207 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP31 VDD net178 net204 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP33 net177 S0 net178 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP22 net184 S0 net198 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP21 VDD C net177 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net184 net201 net183 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 VDD S1 net0188 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP27 net205 S1 net207 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP28 net205 net0188 net204 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD B net183 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP18 VDD A net198 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 VDD D net180 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP17 VDD S0 net201 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP29 VDD net205 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN32 net178 S0 net180 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN30 net207 net184 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN18 net198 A VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN22 net198 net201 net184 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN23 net183 S0 net184 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN21 net177 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN33 net178 net201 net177 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN31 net204 net178 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0188 S1 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN27 net207 net0188 net205 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN28 net204 S1 net205 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN20 net180 D VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN29 Z net205 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 net183 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN17 net201 S0 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends MXB4M2HM
                                                           
.subckt MXB4M4HM Z A B C D S0 S1 VDD VSS 
MP32 net180 net201 net178 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP33 net177 S0 net178 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP30 VDD net184 net207 VDD P_15_LL_EE2_UCFN w=0.71u l=0.12u
MP31 VDD net178 net204 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP22 net184 S0 net198 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP21 VDD C net177 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net184 net201 net183 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP26 VDD S1 net0188 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP27 net205 S1 net207 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP28 net205 net0188 net204 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP19 VDD B net183 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP18 VDD A net198 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP20 VDD D net180 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP17 VDD S0 net201 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP29 VDD net205 Z VDD P_15_LL_EE2_UCFN w=1.34u l=0.12u
MN32 net178 S0 net180 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN30 net207 net184 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN18 net198 A VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN22 net198 net201 net184 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN23 net183 S0 net184 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN21 net177 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN31 net204 net178 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN33 net178 net201 net177 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN26 net0188 S1 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN27 net207 net0188 net205 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN28 net204 S1 net205 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN20 net180 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN29 Z net205 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN19 net183 B VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN17 net201 S0 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
.ends MXB4M4HM
                                                           
.subckt ND2B1M0HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends ND2B1M0HM
                                                           
.subckt ND2B1M12HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 Z B net02 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN2 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=1.15u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=2.91u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.91u l=0.12u
.ends ND2B1M12HM
                                                           
.subckt ND2B1M1HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
.ends ND2B1M1HM
                                                           
.subckt ND2B1M2HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
.ends ND2B1M2HM
                                                           
.subckt ND2B1M4HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z B net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
.ends ND2B1M4HM
                                                           
.subckt ND2B1M8HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
.ends ND2B1M8HM
                                                           
.subckt ND2M0HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends ND2M0HM
                                                           
.subckt ND2M12HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.91u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=2.91u l=0.12u
.ends ND2M12HM
                                                           
.subckt ND2M16HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=3.84u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=3.84u l=0.12u
.ends ND2M16HM
                                                           
.subckt ND2M1HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
.ends ND2M1HM
                                                           
.subckt ND2M2HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
.ends ND2M2HM
                                                           
.subckt ND2M3HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.83u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.83u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.70u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.70u l=0.12u
.ends ND2M3HM
                                                           
.subckt ND2M4HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
.ends ND2M4HM
                                                           
.subckt ND2M5HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.41u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.41u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.22u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.22u l=0.12u
.ends ND2M5HM
                                                           
.subckt ND2M6HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.46u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.46u l=0.12u
.ends ND2M6HM
                                                           
.subckt ND2M8HM Z A B VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
.ends ND2M8HM
                                                           
.subckt ND3B1M0HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z C net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
.ends ND3B1M0HM
                                                           
.subckt ND3B1M1HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 Z C net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends ND3B1M1HM
                                                           
.subckt ND3B1M2HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 B net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z C net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends ND3B1M2HM
                                                           
.subckt ND3B1M4HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 B net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 Z C net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.87u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.87u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.87u l=0.12u
.ends ND3B1M4HM
                                                           
.subckt ND3B1M8HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 B net03 VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MN2 Z C net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=1.96u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.75u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=1.75u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.75u l=0.12u
.ends ND3B1M8HM
                                                           
.subckt ND3M0HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
.ends ND3M0HM
                                                           
.subckt ND3M12HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.62u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=2.62u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=2.62u l=0.12u
.ends ND3M12HM
                                                           
.subckt ND3M16HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=4.38u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=3.50u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=3.50u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=3.50u l=0.12u
.ends ND3M16HM
                                                           
.subckt ND3M1HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends ND3M1HM
                                                           
.subckt ND3M2HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends ND3M2HM
                                                           
.subckt ND3M3HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.85u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
.ends ND3M3HM
                                                           
.subckt ND3M4HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.87u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.87u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.87u l=0.12u
.ends ND3M4HM
                                                           
.subckt ND3M6HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.31u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.31u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=1.31u l=0.12u
.ends ND3M6HM
                                                           
.subckt ND3M8HM Z A B C VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=1.93u l=0.12u
MN2 net02 C VSS VSS N_15_LL_EE2_UCFN w=1.93u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.75u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.75u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=1.75u l=0.12u
.ends ND3M8HM
                                                           
.subckt ND4B1M0HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net03 B net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z D net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends ND4B1M0HM
                                                           
.subckt ND4B1M1HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net03 B net04 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 Z D net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends ND4B1M1HM
                                                           
.subckt ND4B1M2HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net03 B net04 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z D net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends ND4B1M2HM
                                                           
.subckt ND4B1M4HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 B net04 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 Z D net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
.ends ND4B1M4HM
                                                           
.subckt ND4B1M8HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 B net04 VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MN3 Z D net02 VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MN4 net04 net01 VSS VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
.ends ND4B1M8HM
                                                           
.subckt ND4B2M0HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net03 C net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net04 D net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends ND4B2M0HM
                                                           
.subckt ND4B2M1HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net03 C net04 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net04 D net05 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN5 Z net02 net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends ND4B2M1HM
                                                           
.subckt ND4B2M2HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net03 C net04 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net04 D net05 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 Z net02 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends ND4B2M2HM
                                                           
.subckt ND4B2M4HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 C net04 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net04 D net05 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 Z net02 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
.ends ND4B2M4HM
                                                           
.subckt ND4B2M8HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 C net04 VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MN3 net04 D net05 VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MN4 net05 net01 VSS VSS N_15_LL_EE2_UCFN w=2.1u l=0.12u
MN5 Z net02 net03 VSS N_15_LL_EE2_UCFN w=2.1u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
.ends ND4B2M8HM
                                                           
.subckt ND4M0HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends ND4M0HM
                                                           
.subckt ND4M12HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=2.33u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=2.33u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=2.33u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=2.33u l=0.12u
.ends ND4M12HM
                                                           
.subckt ND4M16HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=4.1u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=4.28u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=4.28u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=4.1u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=3.11u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=3.11u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=3.11u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=3.11u l=0.12u
.ends ND4M16HM
                                                           
.subckt ND4M1HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends ND4M1HM
                                                           
.subckt ND4M2HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends ND4M2HM
                                                           
.subckt ND4M4HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=0.78u l=0.12u
.ends ND4M4HM
                                                           
.subckt ND4M6HM Z A B C D VDD VSS 
MN6 net02 C net04 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN4 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net03 net01 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net05 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 A net05 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP6 net02 C VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net06 net02 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net03 net01 net06 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net02 D VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 net01 B VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 net01 A VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 Z net03 VDD VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends ND4M6HM
                                                           
.subckt ND4M8HM Z A B C D VDD VSS 
MN0 Z A net01 VSS N_15_LL_EE2_UCFN w=2.1u l=0.12u
MN1 net01 B net02 VSS N_15_LL_EE2_UCFN w=2.1u l=0.12u
MN2 net02 C net03 VSS N_15_LL_EE2_UCFN w=2.1u l=0.12u
MN3 net03 D VSS VSS N_15_LL_EE2_UCFN w=2.1u l=0.12u
MP0 VDD A Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP1 VDD B Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP2 VDD C Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
MP3 VDD D Z VDD P_15_LL_EE2_UCFN w=1.55u l=0.12u
.ends ND4M8HM
                                                           
.subckt NR2B1M0HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net02 B Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends NR2B1M0HM
                                                           
.subckt NR2B1M12HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=1.17u l=0.12u
MP1 net02 B Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP2 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends NR2B1M12HM
                                                           
.subckt NR2B1M1HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net02 B Z VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP2 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
.ends NR2B1M1HM
                                                           
.subckt NR2B1M2HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net02 B Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR2B1M2HM
                                                           
.subckt NR2B1M4HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 B Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR2B1M4HM
                                                           
.subckt NR2B1M8HM Z B NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 B Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD net01 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends NR2B1M8HM
                                                           
.subckt NR2M0HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends NR2M0HM
                                                           
.subckt NR2M12HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.22u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=2.22u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends NR2M12HM
                                                           
.subckt NR2M16HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.84u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=2.84u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends NR2M16HM
                                                           
.subckt NR2M1HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends NR2M1HM
                                                           
.subckt NR2M2HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR2M2HM
                                                           
.subckt NR2M3HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=1.07u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=1.07u l=0.12u
.ends NR2M3HM
                                                           
.subckt NR2M4HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR2M4HM
                                                           
.subckt NR2M5HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=1.72u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=1.72u l=0.12u
.ends NR2M5HM
                                                           
.subckt NR2M6HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.11u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends NR2M6HM
                                                           
.subckt NR2M8HM Z A B VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1.48u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD B net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends NR2M8HM
                                                           
.subckt NR3B1M0HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net02 C Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends NR3B1M0HM
                                                           
.subckt NR3B1M1HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net02 C Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends NR3B1M1HM
                                                           
.subckt NR3B1M2HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net02 C Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR3B1M2HM
                                                           
.subckt NR3B1M4HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net02 C Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR3B1M4HM
                                                           
.subckt NR3B1M8HM Z B C NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net02 C Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends NR3B1M8HM
                                                           
.subckt NR3M0HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends NR3M0HM
                                                           
.subckt NR3M12HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.88u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1.88u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=1.88u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends NR3M12HM
                                                           
.subckt NR3M16HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2.51u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=2.51u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=2.51u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends NR3M16HM
                                                           
.subckt NR3M1HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends NR3M1HM
                                                           
.subckt NR3M2HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR3M2HM
                                                           
.subckt NR3M4HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR3M4HM
                                                           
.subckt NR3M6HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.94u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends NR3M6HM
                                                           
.subckt NR3M8HM Z A B C VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=1.25u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD C net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends NR3M8HM
                                                           
.subckt NR4B1M0HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net04 B net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 net02 D Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends NR4B1M0HM
                                                           
.subckt NR4B1M1HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 net04 B net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net02 D Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR4B1M1HM
                                                           
.subckt NR4B1M2HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net04 B net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net02 D Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR4B1M2HM
                                                           
.subckt NR4B1M4HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net04 B net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net02 D Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends NR4B1M4HM
                                                           
.subckt NR4B1M8HM Z B C D NA VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net04 B net03 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP3 net02 D Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends NR4B1M8HM
                                                           
.subckt NR4B2M0HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 VDD net01 net05 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP5 net03 net02 Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends NR4B2M0HM
                                                           
.subckt NR4B2M1HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 net03 net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR4B2M1HM
                                                           
.subckt NR4B2M2HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net01 net05 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 net03 net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR4B2M2HM
                                                           
.subckt NR4B2M4HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD net01 net05 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 net03 net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends NR4B2M4HM
                                                           
.subckt NR4B2M8HM Z C D NA NB VDD VSS 
MN0 net01 NA VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 NB VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP0 VDD NA net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD NB net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP4 VDD net01 net05 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP5 net03 net02 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends NR4B2M8HM
                                                           
.subckt NR4M0HM Z A B C D VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 VDD D net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends NR4M0HM
                                                           
.subckt NR4M12HM Z A B C D VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
MP3 VDD D net03 VDD P_15_LL_EE2_UCFN w=8.16u l=0.12u
.ends NR4M12HM
                                                           
.subckt NR4M16HM Z A B C D VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=4u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=4u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=4u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=4u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
MP3 VDD D net03 VDD P_15_LL_EE2_UCFN w=10.88u l=0.12u
.ends NR4M16HM
                                                           
.subckt NR4M1HM Z A B C D VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD D net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends NR4M1HM
                                                           
.subckt NR4M2HM Z A B C D VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD D net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR4M2HM
                                                           
.subckt NR4M4HM Z A B C D VDD VSS 
MN6 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net06 net01 VSS VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN4 net06 net02 net03 VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP6 net01 D net04 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP5 net03 net01 VDD VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 net04 C VDD VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP3 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net05 A VDD VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 net02 B net05 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 Z net03 VDD VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends NR4M4HM
                                                           
.subckt NR4M6HM Z A B C D VDD VSS 
MN6 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net06 net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net06 net02 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP6 net01 D net04 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP5 net03 net01 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net04 C VDD VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP3 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net05 A VDD VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 net02 B net05 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 Z net03 VDD VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends NR4M6HM
                                                           
.subckt NR4M8HM Z A B C D VDD VSS 
MN0 Z A VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN1 Z B VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN2 Z C VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN3 Z D VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP0 net01 A Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP1 net02 B net01 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP2 net03 C net02 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
MP3 VDD D net03 VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends NR4M8HM
                                                           
.subckt OA211M0HM Z A1 A2 B C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA211M0HM
                                                           
.subckt OA211M1HM Z A1 A2 B C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA211M1HM
                                                           
.subckt OA211M2HM Z A1 A2 B C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA211M2HM
                                                           
.subckt OA211M4HM Z A1 A2 B C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA211M4HM
                                                           
.subckt OA211M8HM Z A1 A2 B C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net03 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B net03 VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP3 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP4 VDD net03 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA211M8HM
                                                           
.subckt OA21M0HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA21M0HM
                                                           
.subckt OA21M1HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA21M1HM
                                                           
.subckt OA21M2HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA21M2HM
                                                           
.subckt OA21M4HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA21M4HM
                                                           
.subckt OA21M8HM Z A1 A2 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA21M8HM
                                                           
.subckt OA221M0HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA221M0HM
                                                           
.subckt OA221M1HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA221M1HM
                                                           
.subckt OA221M2HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA221M2HM
                                                           
.subckt OA221M4HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA221M4HM
                                                           
.subckt OA221M8HM Z A1 A2 B1 B2 C VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 Z net03 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP5 VDD net03 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA221M8HM
                                                           
.subckt OA222M0HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 net06 C1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD C2 net06 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA222M0HM
                                                           
.subckt OA222M1HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 net06 C1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD C2 net06 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA222M1HM
                                                           
.subckt OA222M2HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 net06 C1 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD C2 net06 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA222M2HM
                                                           
.subckt OA222M4HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net06 C1 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD C2 net06 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA222M4HM
                                                           
.subckt OA222M8HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 net03 A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net03 A2 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN6 Z net03 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net04 A1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net05 B1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net06 C1 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD C2 net06 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net03 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA222M8HM
                                                           
.subckt OA22M0HM Z A1 A2 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net04 B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA22M0HM
                                                           
.subckt OA22M1HM Z A1 A2 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net04 B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA22M1HM
                                                           
.subckt OA22M2HM Z A1 A2 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net04 B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA22M2HM
                                                           
.subckt OA22M4HM Z A1 A2 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP2 net04 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA22M4HM
                                                           
.subckt OA22M8HM Z A1 A2 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net04 B1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA22M8HM
                                                           
.subckt OA31M0HM Z A1 A2 A3 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA31M0HM
                                                           
.subckt OA31M1HM Z A1 A2 A3 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA31M1HM
                                                           
.subckt OA31M2HM Z A1 A2 A3 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA31M2HM
                                                           
.subckt OA31M4HM Z A1 A2 A3 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.40u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA31M4HM
                                                           
.subckt OA31M8HM Z A1 A2 A3 B VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.92u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.92u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.92u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.92u l=0.12u
MN4 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.80u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA31M8HM
                                                           
.subckt OA32M0HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA32M0HM
                                                           
.subckt OA32M1HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA32M1HM
                                                           
.subckt OA32M2HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA32M2HM
                                                           
.subckt OA32M4HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP4 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=0.60u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA32M4HM
                                                           
.subckt OA32M8HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=1.20u l=0.12u
MP4 VDD B2 net05 VDD P_15_LL_EE2_UCFN w=1.20u l=0.12u
MP5 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA32M8HM
                                                           
.subckt OA33M0HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 net06 B2 net05 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD B3 net06 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OA33M0HM
                                                           
.subckt OA33M1HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 net06 B2 net05 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD B3 net06 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OA33M1HM
                                                           
.subckt OA33M2HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN6 Z net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 net06 B2 net05 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD B3 net06 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP6 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OA33M2HM
                                                           
.subckt OA33M4HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN6 Z net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net06 B2 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD B3 net06 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OA33M4HM
                                                           
.subckt OA33M8HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 net02 A1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net02 A2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 A3 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN6 Z net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net04 A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD A3 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net05 B1 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net06 B2 net05 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD B3 net06 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP6 VDD net02 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OA33M8HM
                                                           
.subckt OAI211B100M0HM Z A1 B C NA2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 Z net01 net03 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
.ends OAI211B100M0HM
                                                           
.subckt OAI211B100M1HM Z A1 B C NA2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN3 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN4 Z net01 net03 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MP0 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OAI211B100M1HM
                                                           
.subckt OAI211B100M2HM Z A1 B C NA2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net03 B net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net02 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net01 net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net04 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI211B100M2HM
                                                           
.subckt OAI211B100M4HM Z A1 B C NA2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN2 net03 B net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net02 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net01 net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net04 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI211B100M4HM
                                                           
.subckt OAI211B100M8HM Z A1 B C NA2 VDD VSS 
MN0 Z A1 net03 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 B net02 VSS N_15_LL_EE2_UCFN w=2.33u l=0.12u
MN3 net02 C VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN4 Z net01 net03 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net04 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
MP4 VDD net01 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OAI211B100M8HM
                                                           
.subckt OAI211M0HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends OAI211M0HM
                                                           
.subckt OAI211M1HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
.ends OAI211M1HM
                                                           
.subckt OAI211M2HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
.ends OAI211M2HM
                                                           
.subckt OAI211M4HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
.ends OAI211M4HM
                                                           
.subckt OAI211M8HM Z A1 A2 B C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net02 B net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net01 C VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
MP3 VDD C Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
.ends OAI211M8HM
                                                           
.subckt OAI21B01M0HM Z A1 A2 NB VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends OAI21B01M0HM
                                                           
.subckt OAI21B01M1HM Z A1 A2 NB VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
.ends OAI21B01M1HM
                                                           
.subckt OAI21B01M2HM Z A1 A2 NB VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
.ends OAI21B01M2HM
                                                           
.subckt OAI21B01M4HM Z A1 A2 NB VDD VSS 
MN0 net02 A1 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net01 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
.ends OAI21B01M4HM
                                                           
.subckt OAI21B01M8HM Z A1 A2 NB VDD VSS 
MN0 net02 A1 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN1 net02 A2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN2 net01 NB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net02 net01 Z VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD NB net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
.ends OAI21B01M8HM
                                                           
.subckt OAI21B10M0HM Z A1 B NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z net01 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
.ends OAI21B10M0HM
                                                           
.subckt OAI21B10M1HM Z A1 B NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 Z net01 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OAI21B10M1HM
                                                           
.subckt OAI21B10M2HM Z A1 B NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 Z net01 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI21B10M2HM
                                                           
.subckt OAI21B10M4HM Z A1 B NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net02 B VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 Z net01 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI21B10M4HM
                                                           
.subckt OAI21B10M8HM Z A1 B NA2 VDD VSS 
MN0 net02 A1 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z B net02 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN3 net02 net01 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
MP3 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OAI21B10M8HM
                                                           
.subckt OAI21B20M0HM Z B NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends OAI21B20M0HM
                                                           
.subckt OAI21B20M1HM Z B NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B net03 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
.ends OAI21B20M1HM
                                                           
.subckt OAI21B20M2HM Z B NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B net03 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
.ends OAI21B20M2HM
                                                           
.subckt OAI21B20M4HM Z B NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z B net03 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
.ends OAI21B20M4HM
                                                           
.subckt OAI21B20M8HM Z B NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z B net03 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
MP3 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
.ends OAI21B20M8HM
                                                           
.subckt OAI21M0HM Z A1 A2 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends OAI21M0HM
                                                           
.subckt OAI21M1HM Z A1 A2 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
.ends OAI21M1HM
                                                           
.subckt OAI21M2HM Z A1 A2 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
.ends OAI21M2HM
                                                           
.subckt OAI21M3HM Z A1 A2 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=1.03u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI21M3HM
                                                           
.subckt OAI21M4HM Z A1 A2 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
.ends OAI21M4HM
                                                           
.subckt OAI21M6HM Z A1 A2 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MN2 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.57u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI21M6HM
                                                           
.subckt OAI21M8HM Z A1 A2 B VDD VSS 
MN0 net01 A1 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN1 net01 A2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN2 Z B net01 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD B Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
.ends OAI21M8HM
                                                           
.subckt OAI221M0HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD C Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends OAI221M0HM
                                                           
.subckt OAI221M1HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD C Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
.ends OAI221M1HM
                                                           
.subckt OAI221M2HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD C Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
.ends OAI221M2HM
                                                           
.subckt OAI221M4HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD C Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
.ends OAI221M4HM
                                                           
.subckt OAI221M8HM Z A1 A2 B1 B2 C VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN4 net01 C VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD C Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
.ends OAI221M8HM
                                                           
.subckt OAI222M0HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP4 net05 C1 Z VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP5 VDD C2 net05 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends OAI222M0HM
                                                           
.subckt OAI222M1HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.40u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 net05 C1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD C2 net05 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OAI222M1HM
                                                           
.subckt OAI222M2HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net05 C1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD C2 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI222M2HM
                                                           
.subckt OAI222M4HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net05 C1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD C2 net05 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI222M4HM
                                                           
.subckt OAI222M8HM Z A1 A2 B1 B2 C1 C2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 Z A2 net02 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net02 B1 net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net02 B2 net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN4 net01 C1 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN5 net01 C2 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD A2 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 net05 C1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 VDD C2 net05 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OAI222M8HM
                                                           
.subckt OAI22B10M0HM Z A1 B1 B2 NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Z net01 net02 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
.ends OAI22B10M0HM
                                                           
.subckt OAI22B10M1HM Z A1 B1 B2 NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN4 Z net01 net02 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OAI22B10M1HM
                                                           
.subckt OAI22B10M2HM Z A1 B1 B2 NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 Z net01 net02 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI22B10M2HM
                                                           
.subckt OAI22B10M4HM Z A1 B1 B2 NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 B1 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 Z net01 net02 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI22B10M4HM
                                                           
.subckt OAI22B10M8HM Z A1 B1 B2 NA2 VDD VSS 
MN0 Z A1 net02 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 B1 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN3 net02 B2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN4 Z net01 net02 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net03 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD NA2 net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD net01 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OAI22B10M8HM
                                                           
.subckt OAI22B20M0HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 Z B2 net03 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends OAI22B20M0HM
                                                           
.subckt OAI22B20M1HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 Z B2 net03 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN4 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
.ends OAI22B20M1HM
                                                           
.subckt OAI22B20M2HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 Z B2 net03 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
.ends OAI22B20M2HM
                                                           
.subckt OAI22B20M4HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 Z B2 net03 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN4 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=0.91u l=0.12u
.ends OAI22B20M4HM
                                                           
.subckt OAI22B20M8HM Z B1 B2 NA1 NA2 VDD VSS 
MN0 net02 NA1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 NA2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 Z B1 net03 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN3 Z B2 net03 VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN4 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 VDD NA1 net02 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP1 VDD NA2 net02 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP2 net04 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 VDD net02 Z VDD P_15_LL_EE2_UCFN w=1.83u l=0.12u
.ends OAI22B20M8HM
                                                           
.subckt OAI22M0HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP2 net03 B1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP3 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
.ends OAI22M0HM
                                                           
.subckt OAI22M1HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net03 B1 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OAI22M1HM
                                                           
.subckt OAI22M2HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net03 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI22M2HM
                                                           
.subckt OAI22M4HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=1.05u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net03 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI22M4HM
                                                           
.subckt OAI22M8HM Z A1 A2 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN2 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MN3 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=2.11u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD A2 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 net03 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B2 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OAI22M8HM
                                                           
.subckt OAI31M0HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 VDD B Z VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends OAI31M0HM
                                                           
.subckt OAI31M1HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD B Z VDD P_15_LL_EE2_UCFN w=0.27u l=0.12u
.ends OAI31M1HM
                                                           
.subckt OAI31M2HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD B Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OAI31M2HM
                                                           
.subckt OAI31M4HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD B Z VDD P_15_LL_EE2_UCFN w=0.76u l=0.12u
.ends OAI31M4HM
                                                           
.subckt OAI31M8HM Z A1 A2 A3 B VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN3 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 VDD B Z VDD P_15_LL_EE2_UCFN w=1.52u l=0.12u
.ends OAI31M8HM
                                                           
.subckt OAI32M0HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
.ends OAI32M0HM
                                                           
.subckt OAI32M1HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP4 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
.ends OAI32M1HM
                                                           
.subckt OAI32M2HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP4 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
.ends OAI32M2HM
                                                           
.subckt OAI32M4HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=1.14u l=0.12u
MP4 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=1.14u l=0.12u
.ends OAI32M4HM
                                                           
.subckt OAI32M8HM Z A1 A2 A3 B1 B2 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP4 VDD B2 net04 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends OAI32M8HM
                                                           
.subckt OAI33M0HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 net05 B2 net04 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP5 VDD B3 net05 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OAI33M0HM
                                                           
.subckt OAI33M1HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 net05 B2 net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP5 VDD B3 net05 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
.ends OAI33M1HM
                                                           
.subckt OAI33M2HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net05 B2 net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD B3 net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OAI33M2HM
                                                           
.subckt OAI33M4HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=0.78u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 net05 B2 net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD B3 net05 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OAI33M4HM
                                                           
.subckt OAI33M8HM Z A1 A2 A3 B1 B2 B3 VDD VSS 
MN0 Z A1 net01 VSS N_15_LL_EE2_UCFN w=1.56u l=0.12u
MN1 Z A2 net01 VSS N_15_LL_EE2_UCFN w=1.64u l=0.12u
MN2 Z A3 net01 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN3 net01 B1 VSS VSS N_15_LL_EE2_UCFN w=1.56u l=0.12u
MN4 net01 B2 VSS VSS N_15_LL_EE2_UCFN w=1.56u l=0.12u
MN5 net01 B3 VSS VSS N_15_LL_EE2_UCFN w=1.56u l=0.12u
MP0 net02 A1 Z VDD P_15_LL_EE2_UCFN w=2.64u l=0.12u
MP1 net03 A2 net02 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP2 VDD A3 net03 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP3 net04 B1 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP4 net05 B2 net04 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 VDD B3 net05 VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OAI33M8HM
                                                           
.subckt OR2M0HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OR2M0HM
                                                           
.subckt OR2M12HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends OR2M12HM
                                                           
.subckt OR2M16HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=4.48u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends OR2M16HM
                                                           
.subckt OR2M1HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OR2M1HM
                                                           
.subckt OR2M2HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OR2M2HM
                                                           
.subckt OR2M4HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OR2M4HM
                                                           
.subckt OR2M6HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.62u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends OR2M6HM
                                                           
.subckt OR2M8HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.74u l=0.12u
MN2 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.16u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OR2M8HM
                                                           
.subckt OR3M0HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OR3M0HM
                                                           
.subckt OR3M12HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.99u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=3.36u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends OR3M12HM
                                                           
.subckt OR3M16HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=4u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends OR3M16HM
                                                           
.subckt OR3M1HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OR3M1HM
                                                           
.subckt OR3M2HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.20u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
.ends OR3M2HM
                                                           
.subckt OR3M4HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OR3M4HM
                                                           
.subckt OR3M6HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends OR3M6HM
                                                           
.subckt OR3M8HM Z A B C VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN3 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OR3M8HM
                                                           
.subckt OR4M0HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
.ends OR4M0HM
                                                           
.subckt OR4M12HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=4.08u l=0.12u
.ends OR4M12HM
                                                           
.subckt OR4M16HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=1.06u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=4u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=5.44u l=0.12u
.ends OR4M16HM
                                                           
.subckt OR4M1HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends OR4M1HM
                                                           
.subckt OR4M2HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends OR4M2HM
                                                           
.subckt OR4M4HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends OR4M4HM
                                                           
.subckt OR4M6HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends OR4M6HM
                                                           
.subckt OR4M8HM Z A B C D VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net01 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Z net01 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 net04 C net03 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP3 VDD D net04 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP4 VDD net01 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends OR4M8HM
                                                           
.subckt OR6M0HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends OR6M0HM
                                                           
.subckt OR6M12HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.9u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=3u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=2.22u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=3u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=3u l=0.12u
.ends OR6M12HM
                                                           
.subckt OR6M1HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
.ends OR6M1HM
                                                           
.subckt OR6M2HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
.ends OR6M2HM
                                                           
.subckt OR6M4HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.97u l=0.12u
.ends OR6M4HM
                                                           
.subckt OR6M6HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=1.21u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.46u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=1.46u l=0.12u
.ends OR6M6HM
                                                           
.subckt OR6M8HM Z A B C D E F VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN1 net01 B VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN2 net01 C VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN3 net04 D VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN4 net04 E VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN5 net04 F VSS VSS N_15_LL_EE2_UCFN w=0.67u l=0.12u
MN6 Z net01 net9 VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN7 net9 net04 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 net02 A net01 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP1 net03 B net02 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP2 VDD C net03 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP3 net05 D net04 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP4 net06 E net05 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP5 VDD F net06 VDD P_15_LL_EE2_UCFN w=1.44u l=0.12u
MP6 VDD net01 Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
MP7 VDD net04 Z VDD P_15_LL_EE2_UCFN w=1.94u l=0.12u
.ends OR6M8HM
                                                           
.subckt SDFCM1HM Q QB CKB D SD SE VDD VSS 
MN17 net11 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net8 CKB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN11 net38 net8 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN9 net38 net42 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN8 VSS net38 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net8 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net44 net11 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN5 net53 D net44 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN4 net50 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN3 net53 SE net50 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN10 net53 net14 net42 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP17 VDD SE net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD CKB net8 VDD P_15_LL_EE2_UCFN w=0.18u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP14 net21 net8 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net21 net14 net38 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP9 VDD net42 net38 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net42 net8 net92 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP3 net93 D net92 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD SE net93 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD SD net102 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net102 net11 net92 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends SDFCM1HM
                                                           
.subckt SDFCM2HM Q QB CKB D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CKB VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN26 net0145 net14 net42 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net0154 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN9 net0154 net42 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 VSS net0154 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net0120 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net0120 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP14 net21 net0120 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net21 net14 net0154 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP26 net42 net0120 net0184 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD net42 net0154 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0154 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends SDFCM2HM
                                                           
.subckt SDFCM4HM Q QB CKB D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 net0120 CKB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN26 net0145 net14 net42 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net0154 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN9 net0154 net42 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 VSS net0154 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net0120 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net0120 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP14 net21 net0120 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net21 net14 net0154 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP26 net42 net0120 net0184 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD net42 net0154 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0154 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends SDFCM4HM
                                                           
.subckt SDFCM8HM Q QB CKB D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN20 net0120 CKB VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN26 net0145 net14 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN11 net0154 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0154 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN8 VSS net0154 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net0120 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP20 VDD CKB net0120 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP14 net21 net0120 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net21 net14 net0154 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP26 net42 net0120 net0184 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD net42 net0154 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0154 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends SDFCM8HM
                                                           
.subckt SDFCQM1HM Q CKB D SD SE VDD VSS 
MN17 net11 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net8 CKB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN11 net38 net8 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN9 net38 net42 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN8 VSS net38 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net8 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net44 net11 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN5 net53 D net44 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN4 net50 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN3 net53 SE net50 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN10 net53 net14 net42 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP17 VDD SE net11 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD CKB net8 VDD P_15_LL_EE2_UCFN w=0.18u l=0.12u
MP14 net21 net8 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net21 net14 net38 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP9 VDD net42 net38 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net42 net8 net92 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP3 net93 D net92 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD SE net93 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD SD net102 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net102 net11 net92 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends SDFCQM1HM
                                                           
.subckt SDFCQM2HM Q CKB D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CKB VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN26 net0145 net14 net42 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net0154 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN9 net0154 net42 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 VSS net0154 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net0120 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net0120 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP14 net21 net0120 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net21 net14 net0154 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP26 net42 net0120 net0184 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD net42 net0154 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0154 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends SDFCQM2HM
                                                           
.subckt SDFCQM4HM Q CKB D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 net0120 CKB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN26 net0145 net14 net42 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net0154 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN9 net0154 net42 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 VSS net0154 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net0120 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net0120 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP14 net21 net0120 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net21 net14 net0154 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP26 net42 net0120 net0184 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD net42 net0154 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0154 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends SDFCQM4HM
                                                           
.subckt SDFCQM8HM Q CKB D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN20 net0120 CKB VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN26 net0145 net14 net42 VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN14 net0171 net14 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN11 net0154 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0154 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN8 VSS net0154 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net0120 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP20 VDD CKB net0120 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP14 net21 net0120 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net21 net14 net0154 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP26 net42 net0120 net0184 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD net42 net0154 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0154 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net14 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends SDFCQM8HM
                                                           
.subckt SDFCQRSM1HM Q CKB D RB SB SD SE VDD VSS 
MP6 VDD net0243 net28 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net28 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 net50 net133 net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD SD net50 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD SE net59 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net59 D net58 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 net113 net130 net58 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD RB net31 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net31 net40 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 VDD net113 net40 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP19 VDD SB net40 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP11 net0243 net127 net40 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD RB net28 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net0243 net130 net22 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net22 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP15 VDD CKB net130 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP23 VDD net28 net22 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP16 VDD net130 net127 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP17 VDD SE net133 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net31 net127 net113 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net94 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net28 RB net88 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net94 net40 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net88 net0243 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net113 net130 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net28 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net22 SB net79 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net115 net127 net113 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net115 SE net118 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN4 net118 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN5 net115 D net124 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN6 net124 net133 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN20 net103 net113 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN19 net40 SB net103 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN11 net40 net130 net0243 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN14 net22 net127 net0243 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net79 net28 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net130 CKB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN16 net127 net130 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net133 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFCQRSM1HM
                                                           
.subckt SDFCQRSM2HM Q CKB D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net49 net62 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net62 net52 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN14 net85 net49 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN11 net94 net52 net20 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net49 net94 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net20 net52 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP26 net62 net52 net131 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net103 net49 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFCQRSM2HM
                                                           
.subckt SDFCQRSM4HM Q CKB D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net49 net62 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net62 net52 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN14 net85 net49 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN11 net94 net52 net20 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net49 net94 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net20 net52 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 net62 net52 net131 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP7 net103 net49 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFCQRSM4HM
                                                           
.subckt SDFCQRSM8HM Q CKB D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN20 net52 CKB VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN26 net68 net49 net62 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.72u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.57u l=0.12u
MN7 net62 net52 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN14 net85 net49 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN11 net94 net52 net20 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP20 VDD CKB net52 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP11 net20 net49 net94 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=1u l=0.12u
MP14 net20 net52 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 net62 net52 net131 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP7 net103 net49 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFCQRSM8HM
                                                           
.subckt SDFCRSM1HM Q QB CKB D RB SB SD SE VDD VSS 
MP6 VDD net0243 net28 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net28 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 net50 net133 net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD SD net50 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD SE net59 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net59 D net58 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 net113 net130 net58 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD RB net31 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net31 net40 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 VDD net113 net40 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP19 VDD SB net40 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP11 net0243 net127 net40 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP9 VDD RB net28 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net0243 net130 net22 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net22 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP18 VDD net22 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP15 VDD CKB net130 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP23 VDD net28 net22 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP16 VDD net130 net127 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP17 VDD SE net133 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 net31 net127 net113 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net94 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net28 RB net88 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net94 net40 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net88 net0243 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net113 net130 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net28 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net22 SB net79 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net115 net127 net113 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net115 SE net118 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN4 net118 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN5 net115 D net124 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN6 net124 net133 VSS VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN20 net103 net113 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN19 net40 SB net103 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN11 net40 net130 net0243 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN14 net22 net127 net0243 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net79 net28 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN18 QB net22 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net130 CKB VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN16 net127 net130 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net133 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFCRSM1HM
                                                           
.subckt SDFCRSM2HM Q QB CKB D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net49 net62 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net62 net52 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN14 net85 net49 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN11 net94 net52 net20 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN18 QB net85 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net49 net94 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net20 net52 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP26 net62 net52 net131 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP18 VDD net85 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP7 net103 net49 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFCRSM2HM
                                                           
.subckt SDFCRSM4HM Q QB CKB D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CKB VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net49 net62 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net62 net52 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN14 net85 net49 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN11 net94 net52 net20 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN18 QB net85 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CKB net52 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net49 net94 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net20 net52 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 net62 net52 net131 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP18 VDD net85 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP7 net103 net49 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFCRSM4HM
                                                           
.subckt SDFCRSM8HM Q QB CKB D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN20 net52 CKB VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN26 net68 net49 net62 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.72u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.57u l=0.12u
MN7 net62 net52 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN14 net85 net49 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN11 net94 net52 net20 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN18 QB net85 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP20 VDD CKB net52 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP11 net20 net49 net94 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.57u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=1u l=0.12u
MP14 net20 net52 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 net62 net52 net131 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP18 VDD net85 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP7 net103 net49 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFCRSM8HM
                                                           
.subckt SDFEM1HM Q QB CK D E SD SE VDD VSS 
MN24 QB net136 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP22 VDD net136 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEM1HM
                                                           
.subckt SDFEM2HM Q QB CK D E SD SE VDD VSS 
MN24 QB net136 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.30u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP22 VDD net136 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEM2HM
                                                           
.subckt SDFEM4HM Q QB CK D E SD SE VDD VSS 
MN24 QB net136 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.30u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP22 VDD net136 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEM4HM
                                                           
.subckt SDFEM8HM Q QB CK D E SD SE VDD VSS 
MN24 QB net136 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.88u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MP22 VDD net136 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=1.1u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends SDFEM8HM
                                                           
.subckt SDFEQM1HM Q CK D E SD SE VDD VSS 
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEQM1HM
                                                           
.subckt SDFEQM2HM Q CK D E SD SE VDD VSS 
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.30u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEQM2HM
                                                           
.subckt SDFEQM4HM Q CK D E SD SE VDD VSS 
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.30u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEQM4HM
                                                           
.subckt SDFEQM8HM Q CK D E SD SE VDD VSS 
MN23 Q net21 VSS VSS N_15_LL_EE2_UCFN w=2.12u l=0.12u
MN22 VSS net136 net9 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN21 net21 net35 net9 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net136 net21 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN19 net25 net32 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net56 net32 net27 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN17 VSS net25 net27 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN16 net25 net56 VSS VSS N_15_LL_EE2_UCFN w=0.88u l=0.12u
MN13 net32 net35 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN12 net35 CK VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN11 net38 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net41 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN9 net44 net41 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN8 net53 SE net44 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN7 net50 net38 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net53 net71 net50 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net56 net35 net53 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN4 net59 E VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN3 net62 net136 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN2 net71 net59 net62 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net68 E VSS VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MN0 net71 D net68 VSS N_15_LL_EE2_UCFN w=0.27u l=0.12u
MP21 VDD net21 Q VDD P_15_LL_EE2_UCFN w=2.86u l=0.12u
MP20 net78 net136 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 net78 net32 net21 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP18 VDD net21 net136 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 net21 net35 net25 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP16 VDD net56 net25 VDD P_15_LL_EE2_UCFN w=1.1u l=0.12u
MP15 net93 net35 net56 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net93 net25 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net35 net32 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD CK net35 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 VDD SE net38 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SD net41 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP9 net119 net32 net56 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP8 net114 net71 net119 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD SE net114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP6 net120 net38 net119 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP5 VDD net41 net120 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP4 VDD E net59 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net129 D net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 net132 E net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP1 VDD net59 net129 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net136 net132 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends SDFEQM8HM
                                                           
.subckt SDFEQRM1HM Q CK D E RB SD SE VDD VSS 
MN21 Q net0120 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN20 net0161 net063 net058 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0161 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN18 net051 RB VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN17 net0120 net058 net051 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN0 net080 net066 net058 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN16 net080 net084 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN12 net063 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net066 net063 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net069 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net072 SE VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN15 net075 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net084 net066 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net075 net080 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net084 net063 net099 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN5 net097 net072 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 net099 SE net0105 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net093 net0161 net097 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net096 E net097 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net099 D net096 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN3 net099 net069 net093 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN7 net0105 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP30 VDD net0120 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP29 net058 net066 net0161 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP28 VDD net0120 net0161 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP27 VDD RB net0120 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP26 VDD net058 net0120 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP0 net058 net063 net080 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP25 VDD net084 net080 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP24 net0135 net063 net084 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0135 net080 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD CK net063 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net063 net066 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD E net069 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 VDD SE net072 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP16 net0151 net072 net23 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP15 VDD SD net0151 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP12 net24 E net23 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP13 net18 D net23 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP11 net27 net0161 net24 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SE net27 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net23 net066 net084 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP14 net27 net069 net18 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFEQRM1HM
                                                           
.subckt SDFEQRM2HM Q CK D E RB SD SE VDD VSS 
MN21 Q net0120 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 net0161 net063 net058 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0161 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN18 net051 RB VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN17 net0120 net058 net051 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net080 net066 net058 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN16 net080 net084 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN12 net063 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net066 net063 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net069 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net072 SE VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN15 net075 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net084 net066 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net075 net080 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net084 net063 net099 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN5 net097 net072 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 net099 SE net0105 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net093 net0161 net097 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net096 E net097 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN1 net099 D net096 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net099 net069 net093 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0105 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP30 VDD net0120 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP29 net058 net066 net0161 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP28 VDD net0120 net0161 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP27 VDD RB net0120 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP26 VDD net058 net0120 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP0 net058 net063 net080 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP25 VDD net084 net080 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP24 net0135 net063 net084 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0135 net080 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD CK net063 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net063 net066 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD E net069 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 VDD SE net072 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP16 net0151 net072 net23 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP15 VDD SD net0151 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP12 net24 E net23 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP13 net18 D net23 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP11 net27 net0161 net24 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SE net27 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net23 net066 net084 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP14 net27 net069 net18 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFEQRM2HM
                                                           
.subckt SDFEQRM4HM Q CK D E RB SD SE VDD VSS 
MN21 Q net0120 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN20 net0161 net063 net058 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0161 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN18 net051 RB VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN17 net0120 net058 net051 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net080 net066 net058 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN16 net080 net084 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN12 net063 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net066 net063 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net069 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net072 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net075 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net084 net066 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net075 net080 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net084 net063 net099 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN5 net097 net072 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN6 net099 SE net0105 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net093 net0161 net097 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net096 E net097 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net099 D net096 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net099 net069 net093 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0105 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP30 VDD net0120 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP29 net058 net066 net0161 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP28 VDD net0120 net0161 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP27 VDD RB net0120 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP26 VDD net058 net0120 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP0 net058 net063 net080 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP25 VDD net084 net080 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP24 net0135 net063 net084 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0135 net080 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD CK net063 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net063 net066 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD E net069 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 VDD SE net072 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 net0151 net072 net23 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP15 VDD SD net0151 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP12 net24 E net23 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP13 net18 D net23 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP11 net27 net0161 net24 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SE net27 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net23 net066 net084 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP14 net27 net069 net18 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFEQRM4HM
                                                           
.subckt SDFEQRM8HM Q CK D E RB SD SE VDD VSS 
MN21 Q net0120 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN20 net0161 net063 net058 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0161 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN18 net051 RB VSS VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
MN17 net0120 net058 net051 VSS N_15_LL_EE2_UCFN w=1.1u l=0.12u
MN0 net080 net066 net058 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN16 net080 net084 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN12 net063 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net066 net063 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN10 net069 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net072 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net075 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net084 net066 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net075 net080 net082 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net084 net063 net099 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN5 net097 net072 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN6 net099 SE net0105 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net093 net0161 net097 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net096 E net097 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net099 D net096 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net099 net069 net093 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0105 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP30 VDD net0120 Q VDD P_15_LL_EE2_UCFN w=2.6u l=0.12u
MP29 net058 net066 net0161 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP28 VDD net0120 net0161 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP27 VDD RB net0120 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP26 VDD net058 net0120 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP0 net058 net063 net080 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP25 VDD net084 net080 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP24 net0135 net063 net084 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0135 net080 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net0135 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD CK net063 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP20 VDD net063 net066 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD E net069 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 VDD SE net072 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 net0151 net072 net23 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP15 VDD SD net0151 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP12 net24 E net23 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP13 net18 D net23 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP11 net27 net0161 net24 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP10 VDD SE net27 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net23 net066 net084 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP14 net27 net069 net18 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFEQRM8HM
                                                           
.subckt SDFEQZRM1HM Q CK D E RB SD SE VDD VSS 
MP22 VDD RB net84 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP0 VDD Q net25 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net96 net28 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net25 E net84 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net28 D net84 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD E net96 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 VDD net114 net37 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP6 net37 net117 net36 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP7 VDD SE net43 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP8 net43 net84 net36 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP9 net36 net123 net99 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP10 VDD SD net114 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 VDD SE net117 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 VDD net120 net123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 net64 net128 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP15 net64 net120 net99 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net99 net128 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP17 net136 net120 net128 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP18 VDD net136 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 net10 net123 net136 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net10 Q VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 VSS RB net88 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net84 D net87 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN1 net87 E net88 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN2 net84 net96 net93 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN3 net93 Q net88 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN4 net96 E VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net99 net120 net102 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN6 net102 net84 net105 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN7 net105 net117 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN8 net102 SE net111 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN9 net111 net114 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN10 net114 SD VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net117 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN13 net123 net120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net128 net99 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN17 VSS net128 net130 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN18 net99 net123 net130 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net128 net123 net136 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN20 Q net136 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net136 net120 net79 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 VSS Q net79 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFEQZRM1HM
                                                           
.subckt SDFEQZRM2HM Q CK D E RB SD SE VDD VSS 
MN25 Q net18 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 net122 net18 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN24 net122 net72 net46 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net18 net46 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 VSS net20 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net24 SE net27 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net27 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN21 net30 net72 net24 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net36 net69 net24 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 net36 net48 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN16 net20 net30 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN18 net30 net75 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net20 net75 net46 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net48 net54 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN26 VSS RB net58 VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN0 net54 D net57 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net57 E net58 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net54 net66 net63 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net63 net122 net58 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net66 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net69 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net72 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN13 net75 net72 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP26 VDD net18 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP24 VDD net18 net122 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 net46 net75 net122 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 VDD net46 net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 net30 net75 net94 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP9 net94 SE net36 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net97 net69 net94 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP7 VDD SD net97 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP6 VDD net48 net36 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP5 VDD net54 net48 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP19 net46 net72 net20 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP17 net112 net72 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net30 net20 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 net112 net20 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net122 net130 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net66 net133 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP2 net130 E net54 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net133 D net54 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP4 VDD E net66 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD SE net69 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net72 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 VDD net72 net75 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEQZRM2HM
                                                           
.subckt SDFEQZRM4HM Q CK D E RB SD SE VDD VSS 
MN25 Q net18 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN23 net122 net18 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN24 net122 net72 net46 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net18 net46 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 VSS net20 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net24 SE net27 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 net27 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN21 net30 net72 net24 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net36 net69 net24 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 net36 net48 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN16 net20 net30 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN18 net30 net75 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net20 net75 net46 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net48 net54 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN26 VSS RB net58 VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN0 net54 D net57 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net57 E net58 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net54 net66 net63 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN3 net63 net122 net58 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN4 net66 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net69 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net72 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN13 net75 net72 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP26 VDD net18 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP24 VDD net18 net122 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 net46 net75 net122 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 VDD net46 net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 net30 net75 net94 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP9 net94 SE net36 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net97 net69 net94 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP7 VDD SD net97 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP6 VDD net48 net36 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP5 VDD net54 net48 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP19 net46 net72 net20 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP17 net112 net72 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net30 net20 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP16 net112 net20 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net122 net130 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net66 net133 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP2 net130 E net54 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP3 net133 D net54 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP4 VDD E net66 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD SE net69 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net72 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 VDD net72 net75 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFEQZRM4HM
                                                           
.subckt SDFEQZRM8HM Q CK D E RB SD SE VDD VSS 
MN25 Q net18 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN23 net122 net18 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN24 net122 net72 net46 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net18 net46 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN20 VSS net20 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net24 SE net27 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN9 net27 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN21 net30 net72 net24 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN7 net36 net69 net24 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN6 net36 net48 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN16 net20 net30 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN18 net30 net75 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net20 net75 net46 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN5 net48 net54 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN26 VSS RB net58 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN0 net54 D net57 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net57 E net58 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN2 net54 net66 net63 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN3 net63 net122 net58 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net66 E VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN15 net69 SE VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN12 net72 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN13 net75 net72 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MP26 VDD net18 Q VDD P_15_LL_EE2_UCFN w=2.8u l=0.12u
MP24 VDD net18 net122 VDD P_15_LL_EE2_UCFN w=0.22u l=0.12u
MP25 net46 net75 net122 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 VDD net46 net18 VDD P_15_LL_EE2_UCFN w=1.4u l=0.12u
MP21 net30 net75 net94 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 net94 SE net36 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP8 net97 net69 net94 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MP7 VDD SD net97 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MP6 VDD net48 net36 VDD P_15_LL_EE2_UCFN w=0.69u l=0.12u
MP5 VDD net54 net48 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP19 net46 net72 net20 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP17 net112 net72 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net30 net20 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP16 net112 net20 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 VDD RB net54 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD net122 net130 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD net66 net133 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 net130 E net54 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net133 D net54 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP4 VDD E net66 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD SE net69 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP12 VDD CK net72 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP13 VDD net72 net75 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends SDFEQZRM8HM
                                                           
.subckt SDFERM1HM Q QB CK D E RB SD SE VDD VSS 
MP1 VDD net21 QB VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP14 net23 net118 net26 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net28 net121 net103 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP10 VDD SE net23 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP11 net23 net21 net29 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net26 D net28 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP12 net29 E net28 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP15 VDD SD net35 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP16 net35 net115 net28 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP18 VDD SE net115 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD E net118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net124 net121 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD CK net124 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 VDD RB net49 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net49 net105 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 net49 net124 net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP25 VDD net103 net105 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net131 net124 net105 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
MP26 VDD net131 net64 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP27 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP28 VDD net64 net21 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP29 net131 net121 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP30 VDD net64 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MN22 QB net21 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN7 net82 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net88 net118 net94 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net88 D net91 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN2 net91 E net92 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net94 net21 net92 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net88 SE net82 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net92 net115 VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN8 net103 net124 net88 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN14 net112 net105 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net103 net121 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net112 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net115 SE VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net118 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net121 net124 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net124 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net105 net103 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net105 net121 net131 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN17 net64 net131 net145 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN19 net21 net64 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net21 net124 net131 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 Q net64 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN18 net145 RB VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFERM1HM
                                                           
.subckt SDFERM2HM Q QB CK D E RB SD SE VDD VSS 
MP1 VDD net21 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net23 net118 net26 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net28 net121 net103 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP10 VDD SE net23 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP11 net23 net21 net29 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net26 D net28 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP12 net29 E net28 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP15 VDD SD net35 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP16 net35 net115 net28 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP18 VDD SE net115 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP19 VDD E net118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net124 net121 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD CK net124 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 VDD RB net49 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net49 net105 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 net49 net124 net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP25 VDD net103 net105 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net131 net124 net105 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 VDD net131 net64 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP27 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP28 VDD net64 net21 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP29 net131 net121 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP30 VDD net64 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN22 QB net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net82 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net88 net118 net94 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net88 D net91 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net91 E net92 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net94 net21 net92 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net88 SE net82 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net92 net115 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net103 net124 net88 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN14 net112 net105 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net103 net121 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net112 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net115 SE VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net118 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net121 net124 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net124 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net105 net103 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net105 net121 net131 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN17 net64 net131 net145 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 net21 net64 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net21 net124 net131 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 Q net64 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN18 net145 RB VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
.ends SDFERM2HM
                                                           
.subckt SDFERM4HM Q QB CK D E RB SD SE VDD VSS 
MP1 VDD net21 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP14 net23 net118 net26 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net28 net121 net103 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP10 VDD SE net23 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP11 net23 net21 net29 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net26 D net28 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP12 net29 E net28 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP15 VDD SD net35 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP16 net35 net115 net28 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP18 VDD SE net115 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD E net118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net124 net121 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD CK net124 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 VDD RB net49 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net49 net105 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 net49 net124 net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP25 VDD net103 net105 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net131 net124 net105 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 VDD net131 net64 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP27 VDD RB net64 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP28 VDD net64 net21 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP29 net131 net121 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP30 VDD net64 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MN22 QB net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net82 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net88 net118 net94 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net88 D net91 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net91 E net92 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net94 net21 net92 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net88 SE net82 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net92 net115 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net103 net124 net88 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN14 net112 net105 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net103 net121 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net112 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net115 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net118 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net121 net124 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net124 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net105 net103 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net105 net121 net131 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN17 net64 net131 net145 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 net21 net64 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net21 net124 net131 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 Q net64 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN18 net145 RB VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
.ends SDFERM4HM
                                                           
.subckt SDFERM8HM Q QB CK D E RB SD SE VDD VSS 
MP1 VDD net21 QB VDD P_15_LL_EE2_UCFN w=2.6u l=0.12u
MP14 net23 net118 net26 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP17 net28 net121 net103 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP10 VDD SE net23 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP11 net23 net21 net29 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP13 net26 D net28 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP12 net29 E net28 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP15 VDD SD net35 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP16 net35 net115 net28 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP18 VDD SE net115 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD E net118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD net124 net121 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD CK net124 VDD P_15_LL_EE2_UCFN w=0.55u l=0.12u
MP22 VDD RB net49 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net49 net105 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 net49 net124 net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP25 VDD net103 net105 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net131 net124 net105 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP26 VDD net131 net64 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP27 VDD RB net64 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP28 VDD net64 net21 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP29 net131 net121 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP30 VDD net64 Q VDD P_15_LL_EE2_UCFN w=2.6u l=0.12u
MN22 QB net21 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN7 net82 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net88 net118 net94 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net88 D net91 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net91 E net92 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net94 net21 net92 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net88 SE net82 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net92 net115 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net103 net124 net88 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN14 net112 net105 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net103 net121 net107 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net112 RB VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN9 net115 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net118 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net121 net124 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 net124 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN16 net105 net103 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net105 net121 net131 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN17 net64 net131 net145 VSS N_15_LL_EE2_UCFN w=1.1u l=0.12u
MN19 net21 net64 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net21 net124 net131 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 Q net64 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN18 net145 RB VSS VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
.ends SDFERM8HM
                                                           
.subckt SDFEZRM1HM Q QB CK D E RB SD SE VDD VSS 
MN22 Q net18 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN23 QB net0438 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 net9 net72 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN15 net0438 net18 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN21 net0438 net36 net22 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net18 net22 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 net26 net33 net22 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN18 net57 net33 net28 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN17 VSS net26 net28 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net26 net57 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN13 net33 net36 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net36 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net39 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net45 SD VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN8 net54 SE net45 VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN7 net51 net39 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN6 net54 net9 net51 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN5 net57 net36 net54 VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN4 net60 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net63 net0438 net70 VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN2 net72 net60 net63 VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN1 net69 E net70 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net72 D net69 VSS N_15_LL_EE2_UCFN w=0.45u l=0.12u
MN26 VSS RB net70 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 VDD net18 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP26 VDD net0438 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP23 VDD net18 net0438 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP21 VDD net72 net9 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP24 net22 net33 net0438 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net22 net18 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP17 net22 net36 net26 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP16 VDD net57 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 net97 net36 net57 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP14 net97 net26 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net36 net33 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net36 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD SE net39 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP8 net115 net9 net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD SE net115 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP6 net121 net39 net120 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP5 VDD SD net121 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP4 VDD E net60 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net130 D net72 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP2 net133 E net72 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net60 net130 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP0 VDD net0438 net133 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP9 net120 net33 net57 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP22 VDD RB net72 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends SDFEZRM1HM
                                                           
.subckt SDFEZRM2HM Q QB CK D E RB SD SE VDD VSS 
MP10 VDD net27 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 VDD net85 net82 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net85 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD SE net109 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD E net88 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net20 D net100 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP2 net23 E net100 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net88 net20 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net27 net23 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP22 VDD RB net100 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP16 net47 net138 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net130 net138 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 net47 net85 net130 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net116 net85 net138 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP5 VDD net100 net112 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 VDD net112 net124 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP7 VDD SD net62 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP8 net62 net109 net65 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP9 net65 SE net124 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP21 net130 net82 net65 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP23 VDD net116 net142 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP25 net116 net82 net27 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 VDD net142 net27 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP26 VDD net142 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN8 QB net27 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net82 net85 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net85 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net109 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net88 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net91 net27 net98 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net100 net88 net91 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net97 E net98 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net100 D net97 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN26 VSS RB net98 VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN5 net112 net100 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN19 net138 net82 net116 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net130 net82 net140 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net138 net130 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net124 net112 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net124 net109 net136 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN21 net130 net85 net136 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net133 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN14 net136 SE net133 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN20 VSS net138 net140 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net142 net116 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN24 net27 net85 net116 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net27 net142 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN25 Q net142 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
.ends SDFEZRM2HM
                                                           
.subckt SDFEZRM4HM Q QB CK D E RB SD SE VDD VSS 
MP10 VDD net27 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 VDD net85 net82 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD CK net85 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD SE net109 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD E net88 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP3 net20 D net100 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP2 net23 E net100 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net88 net20 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net27 net23 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP22 VDD RB net100 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP16 net47 net138 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net130 net138 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP17 net47 net85 net130 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net116 net85 net138 VDD P_15_LL_EE2_UCFN w=0.59u l=0.12u
MP5 VDD net100 net112 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 VDD net112 net124 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP7 VDD SD net62 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP8 net62 net109 net65 VDD P_15_LL_EE2_UCFN w=0.19u l=0.12u
MP9 net65 SE net124 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP21 net130 net82 net65 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP23 VDD net116 net142 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP25 net116 net82 net27 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 VDD net142 net27 VDD P_15_LL_EE2_UCFN w=0.63u l=0.12u
MP26 VDD net142 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MN8 QB net27 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net82 net85 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net85 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net109 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net88 E VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net91 net27 net98 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN2 net100 net88 net91 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN1 net97 E net98 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net100 D net97 VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN26 VSS RB net98 VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN5 net112 net100 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN19 net138 net82 net116 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net130 net82 net140 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net138 net130 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net124 net112 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net124 net109 net136 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN21 net130 net85 net136 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net133 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN14 net136 SE net133 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN20 VSS net138 net140 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net142 net116 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN24 net27 net85 net116 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net27 net142 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN25 Q net142 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
.ends SDFEZRM4HM
                                                           
.subckt SDFEZRM8HM Q QB CK D E RB SD SE VDD VSS 
MP10 VDD net27 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 VDD net85 net82 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP12 VDD CK net85 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP15 VDD SE net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 VDD E net88 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net20 D net100 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP2 net23 E net100 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD net88 net20 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP0 VDD net27 net23 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP22 VDD RB net100 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP16 net47 net138 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP18 VDD net130 net138 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP17 net47 net85 net130 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 net116 net85 net138 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP5 VDD net100 net112 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP6 VDD net112 net124 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP7 VDD SD net62 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MP8 net62 net109 net65 VDD P_15_LL_EE2_UCFN w=0.2u l=0.12u
MP9 net65 SE net124 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP21 net130 net82 net65 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP23 VDD net116 net142 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP25 net116 net82 net27 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 VDD net142 net27 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP26 VDD net142 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MN8 QB net27 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN13 net82 net85 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN12 net85 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN15 net109 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net88 E VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net91 net27 net98 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN2 net100 net88 net91 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN1 net97 E net98 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net100 D net97 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN26 VSS RB net98 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN5 net112 net100 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN19 net138 net82 net116 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net130 net82 net140 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN16 net138 net130 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN6 net124 net112 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net124 net109 net136 VSS N_15_LL_EE2_UCFN w=0.23u l=0.12u
MN21 net130 net85 net136 VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN9 net133 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN14 net136 SE net133 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN20 VSS net138 net140 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net142 net116 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN24 net27 net85 net116 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net27 net142 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN25 Q net142 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
.ends SDFEZRM8HM
                                                           
.subckt SDFM1HM Q QB CK D SD SE VDD VSS 
MN17 net11 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net8 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 net0171 net8 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net38 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN9 net38 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN8 VSS net38 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net44 net11 VSS VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN5 net53 D net44 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net50 SD VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net53 SE net50 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN10 net53 net8 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP17 VDD SE net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD CK net8 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 net21 net14 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP11 net21 net8 net38 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net38 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net8 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net42 net14 net92 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net93 D net92 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD SE net93 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD SD net102 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP5 net102 net11 net92 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
.ends SDFM1HM
                                                           
.subckt SDFM2HM Q QB CK D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 net0171 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net0151 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0151 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 VSS net0151 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP14 net21 net14 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP11 net21 net0120 net0151 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net0151 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0151 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
.ends SDFM2HM
                                                           
.subckt SDFM4HM Q QB CK D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN14 net0171 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net0151 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0151 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 VSS net0151 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP14 net21 net14 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net21 net0120 net0151 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net0151 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0151 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.84u l=0.12u
.ends SDFM4HM
                                                           
.subckt SDFM8HM Q QB CK D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN14 net0171 net0120 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0171 net29 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net0151 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0151 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 VSS net0151 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP18 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP14 net21 net14 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=1.1u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net21 net0120 net0151 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net0151 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0151 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=1.68u l=0.12u
.ends SDFM8HM
                                                           
.subckt SDFMM1HM Q QB CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP25 VDD net0242 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0209 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net0209 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN25 QB net0242 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
.ends SDFMM1HM
                                                           
.subckt SDFMM2HM Q QB CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP25 VDD net0242 QB VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0209 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net0209 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN25 QB net0242 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFMM2HM
                                                           
.subckt SDFMM4HM Q QB CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP25 VDD net0242 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0209 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net0209 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN25 QB net0242 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFMM4HM
                                                           
.subckt SDFMM8HM Q QB CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=3.02u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP25 VDD net0242 QB VDD P_15_LL_EE2_UCFN w=2.6u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0210 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0210 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP2 net0210 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN25 QB net0242 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.66u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFMM8HM
                                                           
.subckt SDFMQM1HM Q CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0209 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net0209 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
.ends SDFMQM1HM
                                                           
.subckt SDFMQM2HM Q CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0209 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net0209 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.17u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFMQM2HM
                                                           
.subckt SDFMQM4HM Q CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0209 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net0209 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFMQM4HM
                                                           
.subckt SDFMQM8HM Q CK D1 D2 S SD SE VDD VSS 
MP26 net086 net0251 net056 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0249 net0248 net0189 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP21 VDD net0127 net0189 VDD P_15_LL_EE2_UCFN w=0.67u l=0.12u
MP19 net0181 net0251 net0249 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 net0181 net0242 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD net0249 Q VDD P_15_LL_EE2_UCFN w=3.02u l=0.12u
MP13 net084 net0127 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP22 net0242 net0249 VDD VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net086 net0127 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP14 net084 net0248 net086 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 VDD S net043 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 VDD SE net049 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD SE net0210 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 net0210 net043 net048 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP6 net048 D1 net056 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net051 net049 net056 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 VDD SD net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP5 net057 S net056 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP4 VDD CK net0248 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net0248 net0251 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP2 net0210 D2 net057 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN21 net0255 net0127 VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN17 Q net0249 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN19 VSS net0242 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net0101 net0248 net086 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN22 VSS net0249 net0242 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 net0255 net0251 net0249 VSS N_15_LL_EE2_UCFN w=0.66u l=0.12u
MN20 net0249 net0248 net0244 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net086 net0251 net0129 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0127 net086 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net043 S VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN10 net049 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN5 net0171 S net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net0101 SE net092 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN6 net080 D2 net075 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net075 net049 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN13 VSS net0127 net0129 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net0101 net043 net080 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net092 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net0248 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN1 net0251 net0248 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net0101 D1 net0171 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFMQM8HM
                                                           
.subckt SDFQM1HM Q CK D SD SE VDD VSS 
MN34 net134 net125 net141 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN35 VSS net158 net141 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN19 net125 net128 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN20 net128 CK VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN21 net131 SE VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN24 net158 net125 net123 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN38 net123 net128 net117 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN39 VSS net113 net117 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN40 net113 net123 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN26 net143 SE net146 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN27 net146 SD VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 net149 net131 VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN28 net143 D net149 VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN37 net134 net128 net155 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN31 net155 net143 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN33 net158 net134 VSS VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN32 Q net123 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP35 net210 net158 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 VDD net128 net125 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP20 VDD CK net128 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP21 VDD SE net131 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP24 net123 net128 net158 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP37 net165 net113 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP38 VDD net123 net113 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP39 net165 net125 net123 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 net192 D net143 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP26 VDD SE net192 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP29 net198 net131 net143 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP28 VDD SD net198 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP33 VDD net134 net158 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP30 VDD net143 net185 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP36 net134 net125 net185 VDD P_15_LL_EE2_UCFN w=0.37u l=0.12u
MP34 net210 net128 net134 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP32 VDD net123 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends SDFQM1HM
                                                           
.subckt SDFQM2HM Q CK D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN32 Q net0117 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN40 net0117 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN39 VSS net0117 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN11 net0102 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0102 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN38 net21 net0120 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 VSS net0102 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP37 net0166 net0117 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP38 VDD net21 net0117 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP39 net0166 net14 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net21 net0120 net0102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net0102 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0102 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP32 VDD net0117 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends SDFQM2HM
                                                           
.subckt SDFQM4HM Q CK D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN32 Q net0117 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN40 net0117 net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN39 VSS net0117 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN11 net0102 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0102 net42 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN38 net21 net0120 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 VSS net0102 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP37 net0166 net0117 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP38 VDD net21 net0117 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP39 net0166 net14 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net21 net0120 net0102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net0102 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0102 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP32 VDD net0117 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends SDFQM4HM
                                                           
.subckt SDFQM8HM Q CK D SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN32 Q net0117 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN40 net0117 net21 VSS VSS N_15_LL_EE2_UCFN w=0.6u l=0.12u
MN39 VSS net0117 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN11 net0102 net14 net21 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN9 net0102 net42 VSS VSS N_15_LL_EE2_UCFN w=0.38u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN38 net21 net0120 net0121 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 VSS net0102 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP37 net0166 net0117 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP38 VDD net21 net0117 VDD P_15_LL_EE2_UCFN w=0.69u l=0.12u
MP39 net0166 net14 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net21 net0120 net0102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP9 VDD net42 net0102 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP8 net84 net0102 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP32 VDD net0117 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends SDFQM8HM
                                                           
.subckt SDFQRM1HM Q CK D RB SD SE VDD VSS 
MN24 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN23 VSS net29 net0240 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0118 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net29 net21 net0111 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN17 net0124 SE VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN15 net8 CK VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN21 net0111 RB VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN11 net0142 net14 net21 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN22 net21 net8 net0240 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net0142 net0164 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 net0118 net0142 net0146 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net0164 net14 net0146 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net0151 net0124 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net0160 D net0151 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net0157 SD VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN3 net0160 SE net0157 VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN10 net0160 net8 net0164 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MP24 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP19 VDD RB net0169 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0297 net14 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 net0297 net29 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD SE net0124 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP15 VDD CK net8 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP21 VDD RB net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP11 net21 net8 net0142 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 VDD net0164 net0142 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP8 net0169 net0142 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0169 net8 net0164 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net0164 net14 net0208 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net0209 D net0208 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP4 VDD SD net0218 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP5 net0218 net0124 net0208 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
.ends SDFQRM1HM
                                                           
.subckt SDFQRM2HM Q CK D RB SD SE VDD VSS 
MN24 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 VSS net29 net0240 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0118 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN20 net29 net21 net0111 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN17 net0124 SE VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN15 net8 CK VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN21 net0111 RB VSS VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN11 net0142 net14 net21 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN22 net21 net8 net0240 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net0142 net0164 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN8 net0118 net0142 net0146 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net0164 net14 net0146 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net0151 net0124 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net0160 D net0151 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net0157 SD VSS VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN3 net0160 SE net0157 VSS N_15_LL_EE2_UCFN w=0.2u l=0.12u
MN10 net0160 net8 net0164 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MP24 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD RB net0169 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP23 net0297 net14 net21 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 net0297 net29 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP17 VDD SE net0124 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP15 VDD CK net8 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP21 VDD RB net29 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP11 net21 net8 net0142 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 VDD net0164 net0142 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP8 net0169 net0142 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0169 net8 net0164 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net0164 net14 net0208 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net0209 D net0208 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD SE net0209 VDD P_15_LL_EE2_UCFN w=0.52u l=0.12u
MP4 VDD SD net0218 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
MP5 net0218 net0124 net0208 VDD P_15_LL_EE2_UCFN w=0.24u l=0.12u
.ends SDFQRM2HM
                                                           
.subckt SDFQRM4HM Q CK D RB SD SE VDD VSS 
MN21 net0123 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net0126 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN11 net0132 net0113 net14 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN31 Q net0188 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN23 VSS net0188 net0109 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN9 net0132 net0145 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN32 net0188 net14 net0131 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN33 net0131 RB VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN34 net14 net0120 net0109 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net0126 net0132 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net0145 net0113 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN27 net0141 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0151 net0120 net0145 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net0151 SE net0159 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net0141 net0123 net0151 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN19 net0113 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN25 net0159 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP21 VDD SE net0123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 VDD RB net0180 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net14 net0120 net0132 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP31 VDD net0188 Q VDD P_15_LL_EE2_UCFN w=1.19u l=0.12u
MP32 net0192 net0113 net14 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP33 VDD net14 net0188 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP9 VDD net0145 net0132 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP34 net0192 net0188 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP35 VDD RB net0188 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP8 net0180 net0132 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0180 net0120 net0145 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net0141 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP23 net0199 net0123 net0205 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0199 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0205 SE net0141 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP26 net0145 net0113 net0205 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP19 VDD net0120 net0113 VDD P_15_LL_EE2_UCFN w=0.3u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
.ends SDFQRM4HM
                                                           
.subckt SDFQRM8HM Q CK D RB SD SE VDD VSS 
MN21 net0123 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net0126 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN11 net0132 net0113 net14 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN31 Q net0188 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN23 VSS net0188 net0109 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net0132 net0145 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN32 net0188 net14 net0131 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN33 net0131 RB VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN34 net14 net0120 net0109 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net0126 net0132 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net0145 net0113 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN27 net0141 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0151 net0120 net0145 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net0151 SE net0159 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net0141 net0123 net0151 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN19 net0113 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN25 net0159 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP21 VDD SE net0123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 VDD RB net0180 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net14 net0120 net0132 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP31 VDD net0188 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP32 net0192 net0113 net14 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP33 VDD net14 net0188 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP9 VDD net0145 net0132 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP34 net0192 net0188 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP35 VDD RB net0188 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP8 net0180 net0132 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0180 net0120 net0145 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net0141 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0199 net0123 net0205 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0199 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0205 SE net0141 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP26 net0145 net0113 net0205 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP19 VDD net0120 net0113 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends SDFQRM8HM
                                                           
.subckt SDFQRSM1HM Q CK D RB SB SD SE VDD VSS 
MP6 VDD net0229 net28 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net28 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 net50 net133 net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD SD net50 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD SE net59 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP3 net59 D net58 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP10 net113 net130 net58 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP1 VDD RB net31 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net31 net40 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 VDD net113 net40 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD SB net40 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP11 net0229 net127 net40 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP9 VDD RB net28 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net0229 net130 net22 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net22 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP15 VDD CK net127 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP23 VDD net28 net22 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP16 VDD net127 net130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD SE net133 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net31 net127 net113 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net94 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net28 RB net88 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net94 net40 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net88 net0229 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net113 net130 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net28 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net22 SB net79 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net115 net127 net113 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net115 SE net118 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net118 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net115 D net124 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 net124 net133 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN20 net103 net113 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN19 net40 SB net103 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net40 net130 net0229 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN14 net22 net127 net0229 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net79 net28 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN15 net127 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net130 net127 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net133 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFQRSM1HM
                                                           
.subckt SDFQRSM2HM Q CK D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net52 net62 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net62 net49 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN14 net85 net52 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net94 net49 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net52 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net52 net94 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net20 net49 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP26 net62 net49 net131 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net103 net52 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFQRSM2HM
                                                           
.subckt SDFQRSM4HM Q CK D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net52 net62 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN7 net62 net49 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN14 net85 net52 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net94 net49 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net52 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net52 net94 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net20 net49 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP26 net62 net49 net131 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net103 net52 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFQRSM4HM
                                                           
.subckt SDFQRSM8HM Q CK D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net52 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN26 net68 net52 net62 VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.84u l=0.12u
MN7 net62 net49 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN14 net85 net52 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN11 net94 net49 net20 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP20 VDD CK net52 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net52 net94 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP14 net20 net49 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP26 net62 net49 net131 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net103 net52 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFQRSM8HM
                                                           
.subckt SDFQRXM2HM Q CK D RB SD SE VDD VSS 
MN21 net0123 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net0126 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN11 net0132 net0113 net14 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN31 Q net0188 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 VSS net0188 net0109 VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN9 net0132 net0145 VSS VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN32 net0188 net14 net0131 VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN33 net0131 RB VSS VSS N_15_LL_EE2_UCFN w=0.51u l=0.12u
MN34 net14 net0120 net0109 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN8 net0126 net0132 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net0145 net0113 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN27 net0141 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0151 net0120 net0145 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net0151 SE net0159 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net0141 net0123 net0151 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net0113 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN25 net0159 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP21 VDD SE net0123 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 VDD RB net0180 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net14 net0120 net0132 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP31 VDD net0188 Q VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP32 net0192 net0113 net14 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP33 VDD net14 net0188 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP9 VDD net0145 net0132 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP34 net0192 net0188 VDD VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP35 VDD RB net0188 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 net0180 net0132 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0180 net0120 net0145 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net0141 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP23 net0199 net0123 net0205 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0199 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0205 SE net0141 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP26 net0145 net0113 net0205 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP19 VDD net0120 net0113 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends SDFQRXM2HM
                                                           
.subckt SDFQSM1HM Q CK D SB SD SE VDD VSS 
MN17 net11 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN15 net8 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net0112 net29 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net0171 net8 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net38 net14 net21 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN19 net38 SB net0145 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN20 net0145 net42 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 VSS net38 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net44 net11 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net53 D net44 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net50 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net53 SE net50 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net53 net8 net42 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN21 net0171 SB net0112 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP17 VDD SE net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP23 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP15 VDD CK net8 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP21 VDD SB net0171 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP14 net21 net14 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net21 net8 net38 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP19 VDD SB net38 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP20 VDD net42 net38 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net84 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net8 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net42 net14 net92 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP3 net93 D net92 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP2 VDD SE net93 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD SD net102 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net102 net11 net92 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends SDFQSM1HM
                                                           
.subckt SDFQSM2HM Q CK D SB SD SE VDD VSS 
MP26 net72 net102 net52 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net87 net30 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP1 VDD SB net30 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP24 net52 SE net117 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP22 VDD SD net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP23 net58 net120 net52 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP14 net85 net102 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net117 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net99 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD net99 net102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD net85 net87 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net85 net99 net21 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD SB net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 VDD net72 net21 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 net13 net21 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net13 net99 net72 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD net87 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN0 net93 net87 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net30 net99 net85 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net87 net85 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net21 net102 net85 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 net21 SB net78 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net78 net72 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 VSS net21 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net72 net102 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net30 SB net93 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 Q net87 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN25 net105 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net117 net120 net109 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN24 net109 SE net105 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN26 net109 net99 net72 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN27 net117 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net120 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net99 CK VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN19 net102 net99 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends SDFQSM2HM
                                                           
.subckt SDFQSM4HM Q CK D SB SD SE VDD VSS 
MP26 net72 net102 net52 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net87 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD SB net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 net52 SE net117 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP22 VDD SD net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP23 net58 net120 net52 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP14 net85 net102 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net117 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net99 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD net99 net102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD net85 net87 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net85 net99 net21 VDD P_15_LL_EE2_UCFN w=0.44u l=0.12u
MP2 VDD SB net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 VDD net72 net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net13 net21 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net13 net99 net72 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD net87 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MN0 net93 net87 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net30 net99 net85 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net87 net85 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net21 net102 net85 VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN1 net21 SB net78 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net78 net72 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 VSS net21 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net72 net102 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net30 SB net93 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 Q net87 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN25 net105 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net117 net120 net109 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN24 net109 SE net105 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN26 net109 net99 net72 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN27 net117 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net120 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net99 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net102 net99 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends SDFQSM4HM
                                                           
.subckt SDFQSM8HM Q CK D SB SD SE VDD VSS 
MP26 net72 net102 net52 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net87 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP1 VDD SB net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP24 net52 SE net117 VDD P_15_LL_EE2_UCFN w=0.43u l=0.12u
MP22 VDD SD net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP23 net58 net120 net52 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP14 net85 net102 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net117 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net99 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP19 VDD net99 net102 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net85 net87 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net85 net99 net21 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP2 VDD SB net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 VDD net72 net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net13 net21 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net13 net99 net72 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD net87 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MN0 net93 net87 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN14 net30 net99 net85 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net87 net85 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net21 net102 net85 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net21 SB net78 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net78 net72 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 VSS net21 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net72 net102 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net30 SB net93 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN4 Q net87 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN25 net105 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net117 net120 net109 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN24 net109 SE net105 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN26 net109 net99 net72 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN27 net117 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net120 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net99 CK VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN19 net102 net99 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
.ends SDFQSM8HM
                                                           
.subckt SDFQZRM1HM Q CK D RB SD SE VDD VSS 
MN20 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
.ends SDFQZRM1HM
                                                           
.subckt SDFQZRM2HM Q CK D RB SD SE VDD VSS 
MN24 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends SDFQZRM2HM
                                                           
.subckt SDFQZRM4HM Q CK D RB SD SE VDD VSS 
MN24 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends SDFQZRM4HM
                                                           
.subckt SDFQZRM8HM Q CK D RB SD SE VDD VSS 
MN24 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.91u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.77u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=1.29u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
.ends SDFQZRM8HM
                                                           
.subckt SDFRM1HM Q QB CK D RB SD SE VDD VSS 
MN24 net0174 net29 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net0174 net8 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net0129 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN27 QB net0174 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN20 net29 net21 net0111 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN17 net11 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 net8 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN26 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN21 net0111 RB VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN11 net38 net14 net21 VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN9 net38 net42 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net0129 net38 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net44 net11 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net53 D net44 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net50 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN3 net53 SE net50 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net53 net8 net42 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MP24 VDD net29 net0174 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP25 net21 net14 net0174 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP19 VDD RB net84 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD net0174 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP20 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP17 VDD SE net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP15 VDD CK net8 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP26 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP21 VDD RB net29 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP11 net21 net8 net38 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP9 VDD net42 net38 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP8 net84 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net8 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net42 net14 net92 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP3 net93 D net92 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP2 VDD SE net93 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD SD net102 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net102 net11 net92 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
.ends SDFRM1HM
                                                           
.subckt SDFRM2HM Q QB CK D RB SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net0153 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 net0207 net0142 net0147 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN18 QB net0201 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN30 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN14 net0201 net0120 net0142 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0201 net0207 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN11 net0138 net14 net0142 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN9 net0138 net42 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net0153 net0138 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net0207 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 VDD RB net0210 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP29 VDD net0142 net0207 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP18 VDD net0201 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP30 VDD RB net0207 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net0142 net14 net0201 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net0207 net0201 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 net0142 net0120 net0138 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP9 VDD net42 net0138 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net0210 net0138 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0210 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net0207 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFRM2HM
                                                           
.subckt SDFRM4HM Q QB CK D RB SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net0153 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 net0207 net0142 net0147 VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN18 QB net0201 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN30 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=1.08u l=0.12u
MN14 net0201 net0120 net0142 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0201 net0207 VSS VSS N_15_LL_EE2_UCFN w=0.41u l=0.12u
MN11 net0138 net14 net0142 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN9 net0138 net42 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net0153 net0138 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net0207 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 VDD RB net0210 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP29 VDD net0142 net0207 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP18 VDD net0201 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP30 VDD RB net0207 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP14 net0142 net14 net0201 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net0207 net0201 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP11 net0142 net0120 net0138 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP9 VDD net42 net0138 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP8 net0210 net0138 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0210 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net0207 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFRM4HM
                                                           
.subckt SDFRM8HM Q QB CK D RB SD SE VDD VSS 
MN19 net14 net0120 VSS VSS N_15_LL_EE2_UCFN w=0.55u l=0.12u
MN20 net0120 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net0114 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN28 net0153 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN29 net0207 net0142 net0147 VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN18 QB net0201 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN30 net0147 RB VSS VSS N_15_LL_EE2_UCFN w=1.04u l=0.12u
MN14 net0201 net0120 net0142 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN13 net0201 net0207 VSS VSS N_15_LL_EE2_UCFN w=0.90u l=0.12u
MN11 net0138 net14 net0142 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN9 net0138 net42 VSS VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN8 net0153 net0138 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net0136 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net0207 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN27 net0111 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net0145 net0120 net42 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net0145 SE net0150 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net0111 net0114 net0145 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net0150 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP19 VDD net0120 net14 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP20 VDD CK net0120 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net0114 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP28 VDD RB net0210 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP29 VDD net0142 net0207 VDD P_15_LL_EE2_UCFN w=1.08u l=0.12u
MP18 VDD net0201 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP30 VDD RB net0207 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP14 net0142 net14 net0201 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP13 VDD net0207 net0201 VDD P_15_LL_EE2_UCFN w=1.10u l=0.12u
MP11 net0142 net0120 net0138 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP9 VDD net42 net0138 VDD P_15_LL_EE2_UCFN w=0.5u l=0.12u
MP8 net0210 net0138 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net0210 net0120 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP0 VDD net0207 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP27 VDD D net0111 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 net0169 net0114 net0184 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net0169 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net0184 SE net0111 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP26 net42 net14 net0184 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
.ends SDFRM8HM
                                                           
.subckt SDFRSM1HM Q QB CK D RB SB SD SE VDD VSS 
MP6 VDD net0240 net28 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net28 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 net50 net133 net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD SD net50 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD SE net59 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP3 net59 D net58 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP10 net113 net130 net58 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP1 VDD RB net31 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net31 net40 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP20 VDD net113 net40 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD SB net40 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP11 net0240 net127 net40 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP9 VDD RB net28 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net0240 net130 net22 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP21 VDD SB net22 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP18 VDD net22 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP15 VDD CK net127 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP23 VDD net28 net22 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP16 VDD net127 net130 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP17 VDD SE net133 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 net31 net127 net113 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MN1 net94 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net28 RB net88 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN8 net94 net40 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net88 net0240 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net113 net130 net98 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net28 VSS VSS N_15_LL_EE2_UCFN w=0.53u l=0.12u
MN21 net22 SB net79 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN10 net115 net127 net113 VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN3 net115 SE net118 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN4 net118 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN5 net115 D net124 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN6 net124 net133 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN20 net103 net113 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN19 net40 SB net103 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net40 net130 net0240 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN14 net22 net127 net0240 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN22 net79 net28 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN18 QB net22 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN15 net127 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net130 net127 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net133 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends SDFRSM1HM
                                                           
.subckt SDFRSM2HM Q QB CK D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net52 net62 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net62 net49 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN14 net85 net52 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net94 net49 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN18 QB net85 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net52 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net52 net94 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net20 net49 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP26 net62 net49 net131 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP18 VDD net85 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP7 net103 net52 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFRSM2HM
                                                           
.subckt SDFRSM4HM Q QB CK D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net52 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net52 net62 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net62 net49 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN14 net85 net52 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net94 net49 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN18 QB net85 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net52 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net52 net94 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP14 net20 net49 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP26 net62 net49 net131 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP18 VDD net85 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP7 net103 net52 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFRSM4HM
                                                           
.subckt SDFRSM8HM Q QB CK D RB SB SD SE VDD VSS 
MN19 net49 net52 VSS VSS N_15_LL_EE2_UCFN w=0.54u l=0.12u
MN20 net52 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net55 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net58 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN26 net68 net52 net62 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN24 net68 SE net70 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net58 net55 net68 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN25 net70 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN1 net46 RB VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN2 net109 RB net37 VSS N_15_LL_EE2_UCFN w=0.93u l=0.12u
MN8 net46 net94 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN9 net37 net20 VSS VSS N_15_LL_EE2_UCFN w=0.93u l=0.12u
MN7 net62 net49 net41 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN0 Q net109 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN3 net85 SB net13 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net25 net62 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN14 net85 net52 net20 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN5 net94 SB net25 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN11 net94 net49 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net13 net109 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN18 QB net85 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP6 VDD net20 net109 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP0 VDD net109 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD RB net103 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net103 net94 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP2 VDD net62 net94 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP3 VDD SB net94 VDD P_15_LL_EE2_UCFN w=0.4u l=0.12u
MP19 VDD net52 net49 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP20 VDD CK net52 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net55 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 VDD D net58 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net20 net52 net94 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net125 net55 net131 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP22 VDD SD net125 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP24 net131 SE net58 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP9 VDD RB net109 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP14 net20 net49 net85 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD SB net85 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP26 net62 net49 net131 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP18 VDD net85 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP5 VDD net109 net85 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP7 net103 net52 net62 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
.ends SDFRSM8HM
                                                           
.subckt SDFSM1HM Q QB CK D SB SD SE VDD VSS 
MN23 QB net0171 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN17 net11 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN16 net14 net8 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN15 net8 CK VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net0112 net29 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN14 net0171 net8 net21 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net29 net21 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net38 net14 net21 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN19 net38 SB net0145 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN20 net0145 net42 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 VSS net38 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net42 net14 net33 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN6 net44 net11 VSS VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net53 D net44 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN4 net50 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN3 net53 SE net50 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN10 net53 net8 net42 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN21 net0171 SB net0112 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 Q net29 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP24 VDD net0171 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP17 VDD SE net11 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP16 VDD net8 net14 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP23 VDD net29 net0171 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP15 VDD CK net8 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP21 VDD SB net0171 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP14 net21 net14 net0171 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP12 VDD net21 net29 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net21 net8 net38 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP19 VDD SB net38 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP20 VDD net42 net38 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 net84 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net84 net8 net42 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net42 net14 net92 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP3 net93 D net92 VDD P_15_LL_EE2_UCFN w=0.45u l=0.12u
MP2 VDD SE net93 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP4 VDD SD net102 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net102 net11 net92 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD net29 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends SDFSM1HM
                                                           
.subckt SDFSM2HM Q QB CK D SB SD SE VDD VSS 
MP26 net72 net102 net52 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net87 net30 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP18 VDD net30 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD SB net30 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP24 net52 SE net117 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP22 VDD SD net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP23 net58 net120 net52 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP14 net85 net102 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net117 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net99 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD net99 net102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD net85 net87 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP11 net85 net99 net21 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD SB net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 VDD net72 net21 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 net13 net21 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net13 net99 net72 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD net87 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MN18 QB net30 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net93 net87 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN14 net30 net99 net85 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net87 net85 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN11 net21 net102 net85 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net21 SB net78 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net78 net72 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 VSS net21 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net72 net102 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net30 SB net93 VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 Q net87 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN25 net105 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net117 net120 net109 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN24 net109 SE net105 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN26 net109 net99 net72 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN27 net117 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net120 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net99 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net102 net99 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends SDFSM2HM
                                                           
.subckt SDFSM4HM Q QB CK D SB SD SE VDD VSS 
MP26 net72 net102 net52 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP0 VDD net87 net30 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP18 VDD net30 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD SB net30 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP24 net52 SE net117 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP22 VDD SD net58 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP23 net58 net120 net52 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP14 net85 net102 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net117 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP21 VDD SE net120 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD CK net99 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 VDD net99 net102 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP12 VDD net85 net87 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP11 net85 net99 net21 VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP2 VDD SB net21 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP3 VDD net72 net21 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP8 net13 net21 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net13 net99 net72 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD net87 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MN18 QB net30 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN0 net93 net87 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 net30 net99 net85 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net87 net85 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN11 net21 net102 net85 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net21 SB net78 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net78 net72 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 VSS net21 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net72 net102 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net30 SB net93 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 Q net87 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN25 net105 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net117 net120 net109 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN24 net109 SE net105 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN26 net109 net99 net72 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN27 net117 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN21 net120 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net99 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN19 net102 net99 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends SDFSM4HM
                                                           
.subckt SDFSM8HM Q QB CK D SB SD SE VDD VSS 
MP26 net72 net102 net52 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP0 VDD net87 net30 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP18 VDD net30 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP1 VDD SB net30 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP24 net52 SE net117 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP22 VDD SD net58 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP23 net58 net120 net52 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP14 net85 net102 net30 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP27 VDD D net117 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP21 VDD SE net120 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP20 VDD CK net99 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP19 VDD net99 net102 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net85 net87 VDD P_15_LL_EE2_UCFN w=1.4u l=0.12u
MP11 net85 net99 net21 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD SB net21 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP3 VDD net72 net21 VDD P_15_LL_EE2_UCFN w=0.53u l=0.12u
MP8 net13 net21 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 net13 net99 net72 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP4 VDD net87 Q VDD P_15_LL_EE2_UCFN w=2.8u l=0.12u
MN18 QB net30 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN0 net93 net87 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN14 net30 net99 net85 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN12 net87 net85 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN11 net21 net102 net85 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN1 net21 SB net78 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN2 net78 net72 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN8 VSS net21 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net72 net102 net76 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN3 net30 SB net93 VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN4 Q net87 VSS VSS N_15_LL_EE2_UCFN w=2u l=0.12u
MN25 net105 SD VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN22 net117 net120 net109 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN24 net109 SE net105 VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN26 net109 net99 net72 VSS N_15_LL_EE2_UCFN w=0.43u l=0.12u
MN27 net117 D VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN21 net120 SE VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN20 net99 CK VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN19 net102 net99 VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
.ends SDFSM8HM
                                                           
.subckt SDFZRM1HM Q QB CK D RB SD SE VDD VSS 
MN20 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN21 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN14 QB net38 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP14 VDD net38 QB VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.21u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
.ends SDFZRM1HM
                                                           
.subckt SDFZRM2HM Q QB CK D RB SD SE VDD VSS 
MN24 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN14 QB net38 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP14 VDD net38 QB VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends SDFZRM2HM
                                                           
.subckt SDFZRM4HM Q QB CK D RB SD SE VDD VSS 
MN24 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN14 QB net38 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP14 VDD net38 QB VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=0.50u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.51u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends SDFZRM4HM
                                                           
.subckt SDFZRM8HM Q QB CK D RB SD SE VDD VSS 
MN24 net48 net23 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN25 net116 net26 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN19 net8 SE VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net17 SD VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN17 net20 SE net17 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN16 net26 net23 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN15 Q net48 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN14 QB net38 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MN13 net38 net48 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN22 VSS net38 net44 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN23 VSS net56 net50 VSS N_15_LL_EE2_UCFN w=0.16u l=0.12u
MN10 net56 net26 net48 VSS N_15_LL_EE2_UCFN w=0.91u l=0.12u
MN7 net56 net116 VSS VSS N_15_LL_EE2_UCFN w=0.77u l=0.12u
MN6 net116 net23 net62 VSS N_15_LL_EE2_UCFN w=0.47u l=0.12u
MN5 net62 net20 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net71 net8 net20 VSS N_15_LL_EE2_UCFN w=0.49u l=0.12u
MN2 net71 RB net14 VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net14 D VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net23 CK VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP19 VDD SE net8 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net75 net8 net20 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP17 VDD SD net75 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP16 VDD net23 net26 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP15 VDD net48 Q VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP14 VDD net38 QB VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
MP13 VDD net48 net38 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 net102 net38 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP11 net102 net26 net48 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP10 net48 net23 net56 VDD P_15_LL_EE2_UCFN w=1.29u l=0.12u
MP9 net108 net23 net116 VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP8 net108 net56 VDD VDD P_15_LL_EE2_UCFN w=0.16u l=0.12u
MP7 VDD net116 net56 VDD P_15_LL_EE2_UCFN w=1.04u l=0.12u
MP6 net62 net26 net116 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP5 VDD net20 net62 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP4 net20 SE net71 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP3 VDD RB net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD D net71 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD CK net23 VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
.ends SDFZRM8HM
                                                           
.subckt TIE0HM Z VDD VSS 
MN0 Z net2 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD net2 net2 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends TIE0HM
                                                           
.subckt TIE1HM Z VDD VSS 
MN0 net2 net2 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD net2 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends TIE1HM
                                                           
.subckt WT2HM VDD VSS
.ends WT2HM

.subckt WTBB2HM VDD VSS VBN VBP
.ends WTBB2HM

.subckt WTBN2HM VDD VSS VBN
.ends WTBN2HM

.subckt WTBP2HM VDD VSS VBP
.ends WTBP2HM
                                                           
.subckt XNR2M0HM Z A B VDD VSS 
MN4 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN3 net03 net01 Z VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN2 net02 A Z VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN1 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN0 net02 net03 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 net03 B VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP3 net02 net01 Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 net03 A Z VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP1 net01 A VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 net02 net03 VDD VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends XNR2M0HM
                                                           
.subckt XNR2M1HM Z A B VDD VSS 
MN4 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN3 net03 net01 Z VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 A Z VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN1 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net02 net03 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP4 net03 B VDD VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP3 net02 net01 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 net03 A Z VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP1 net01 A VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP0 net02 net03 VDD VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends XNR2M1HM
                                                           
.subckt XNR2M2HM Z A B VDD VSS 
MN4 net03 B VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN3 net03 net01 Z VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net02 A Z VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net02 net03 VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MP4 net03 B VDD VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP3 net02 net01 Z VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP2 net03 A Z VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
MP1 net01 A VDD VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP0 net02 net03 VDD VDD P_15_LL_EE2_UCFN w=0.66u l=0.12u
.ends XNR2M2HM
                                                           
.subckt XNR2M4HM Z A B VDD VSS 
MP6 VDD A net052 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD net055 net049 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP4 VDD net21 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP5 VDD B net055 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP8 net21 net052 net055 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 net21 A net049 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MN4 Z net21 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN7 net049 net055 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net052 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net055 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN8 net055 A net21 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net049 net052 net21 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
.ends XNR2M4HM
                                                           
.subckt XNR3M0HM Z A B C VDD VSS 
MN3 net138 B net130 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net123 net130 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net130 net141 net121 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net123 C net121 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net138 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net135 net126 net130 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN1 net135 net138 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN8 net141 C VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 Z net121 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN4 net126 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP5 VDD net130 net123 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP6 net121 C net130 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP4 VDD B net126 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP7 net121 net141 net123 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP3 net130 net126 net138 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP8 VDD C net141 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD A net138 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP2 net130 B net135 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP9 VDD net121 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP1 VDD net138 net135 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
.ends XNR3M0HM
                                                           
.subckt XNR3M1HM Z A B C VDD VSS 
MN3 net138 B net130 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 net123 net130 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net130 net141 net121 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN7 net123 C net121 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN0 net138 A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net135 net126 net130 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN1 net135 net138 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN8 net141 C VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 Z net121 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN4 net126 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP5 VDD net130 net123 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP6 net121 C net130 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 VDD B net126 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP7 net121 net141 net123 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP3 net130 net126 net138 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP8 VDD C net141 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD A net138 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 net130 B net135 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP9 VDD net121 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP1 VDD net138 net135 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
.ends XNR3M1HM
                                                           
.subckt XNR3M2HM Z A B C VDD VSS 
MN3 net138 B net130 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN5 net123 net130 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net130 net141 net121 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN7 net123 C net121 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN0 net138 A VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN2 net135 net126 net130 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net135 net138 VSS VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN8 net141 C VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN9 Z net121 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN4 net126 B VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 VDD net130 net123 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net121 C net130 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP4 VDD B net126 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP7 net121 net141 net123 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 net130 net126 net138 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP8 VDD C net141 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP0 VDD A net138 VDD P_15_LL_EE2_UCFN w=0.61u l=0.12u
MP2 net130 B net135 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP9 VDD net121 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD net138 net135 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends XNR3M2HM
                                                           
.subckt XNR3M4HM Z A B C VDD VSS 
MN3 net138 B net130 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN5 net123 net130 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN6 net130 net141 net121 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN7 net123 C net121 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN0 net138 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net135 net126 net130 VSS N_15_LL_EE2_UCFN w=0.34u l=0.12u
MN1 net135 net138 VSS VSS N_15_LL_EE2_UCFN w=0.44u l=0.12u
MN8 net141 C VSS VSS N_15_LL_EE2_UCFN w=0.25u l=0.12u
MN9 Z net121 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN4 net126 B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MP5 VDD net130 net123 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP6 net121 C net130 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP4 VDD B net126 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP7 net121 net141 net123 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP3 net130 net126 net138 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP8 VDD C net141 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP0 VDD A net138 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 net130 B net135 VDD P_15_LL_EE2_UCFN w=0.41u l=0.12u
MP9 VDD net121 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP1 VDD net138 net135 VDD P_15_LL_EE2_UCFN w=0.54u l=0.12u
.ends XNR3M4HM
                                                           
.subckt XNR4M0HM Z A B C D VDD VSS 
MN14 Z net0148 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN12 net083 net025 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN13 net080 net079 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN9 net0148 net079 net051 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN11 net083 D net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net051 net081 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 net0148 net080 net081 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN10 net025 net022 net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net081 A net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 VSS net041 net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net081 net2 net041 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net022 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net025 C VSS VSS N_15_LL_EE2_UCFN w=0.22u l=0.12u
MN1 net041 B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net2 A VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP14 VDD net0148 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP12 VDD net025 net083 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP11 net079 net022 net083 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP10 net079 D net025 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP13 VDD net079 net080 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP8 net081 net079 net0148 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 net051 net080 net0148 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP7 VDD net081 net051 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP6 net035 net2 net081 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net035 net041 VDD VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 net041 A net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD D net022 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD C net025 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 VDD B net041 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP0 VDD A net2 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends XNR4M0HM
                                                           
.subckt XNR4M1HM Z A B C D VDD VSS 
MN14 Z net0148 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN12 net083 net025 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN13 net080 net079 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net0148 net079 net051 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN11 net083 D net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net051 net081 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net0148 net080 net081 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN10 net025 net022 net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net081 A net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 VSS net041 net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net081 net2 net041 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net022 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net025 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net041 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN0 net2 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP14 VDD net0148 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP12 VDD net025 net083 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP11 net079 net022 net083 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP10 net079 D net025 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP13 VDD net079 net080 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net081 net079 net0148 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP9 net051 net080 net0148 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP7 VDD net081 net051 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP6 net035 net2 net081 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net035 net041 VDD VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 net041 A net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD D net022 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD C net025 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 VDD B net041 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP0 VDD A net2 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends XNR4M1HM
                                                           
.subckt XNR4M2HM Z A B C D VDD VSS 
MN14 Z net0148 VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN12 net083 net025 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN13 net080 net079 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN9 net0148 net079 net051 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN11 net083 D net079 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN7 net051 net081 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN8 net0148 net080 net081 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN10 net025 net022 net079 VSS N_15_LL_EE2_UCFN w=0.36u l=0.12u
MN6 net081 A net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 VSS net041 net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN4 net081 net2 net041 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net022 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net025 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net041 B VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN0 net2 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP14 VDD net0148 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net025 net083 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP11 net079 net022 net083 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP10 net079 D net025 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP13 VDD net079 net080 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP8 net081 net079 net0148 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP9 net051 net080 net0148 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP7 VDD net081 net051 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP6 net035 net2 net081 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP5 net035 net041 VDD VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 net041 A net081 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD D net022 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD C net025 VDD P_15_LL_EE2_UCFN w=0.71u l=0.12u
MP1 VDD B net041 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP0 VDD A net2 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
.ends XNR4M2HM
                                                           
.subckt XNR4M4HM Z A B C D VDD VSS 
MN14 Z net79 VSS VSS N_15_LL_EE2_UCFN w=0.96u l=0.12u
MN13 net0117 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN12 net13 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net16 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN16 net70 D net22 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net22 net16 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN15 net70 net0117 net16 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0138 net70 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN17 net79 net70 net37 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net79 net0138 net47 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net37 net47 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN3 net43 A net47 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net43 net49 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN1 net49 net13 net47 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net49 B VSS VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MP14 VDD net79 Z VDD P_15_LL_EE2_UCFN w=1.46u l=0.12u
MP13 VDD D net0117 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP12 VDD A net13 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP11 VDD C net16 VDD P_15_LL_EE2_UCFN w=0.71u l=0.12u
MP16 net22 net0117 net70 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP9 VDD net16 net22 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP15 net16 D net70 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP7 VDD net70 net0138 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP17 net37 net0138 net79 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP18 net47 net70 net79 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP4 VDD net47 net37 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP3 net47 net13 net43 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP2 VDD net49 net43 VDD P_15_LL_EE2_UCFN w=0.31u l=0.12u
MP1 net47 A net49 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP0 VDD B net49 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
.ends XNR4M4HM
                                                           
.subckt XOR2M0HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
.ends XOR2M0HM
                                                           
.subckt XOR2M1HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
.ends XOR2M1HM
                                                           
.subckt XOR2M2HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
.ends XOR2M2HM
                                                           
.subckt XOR2M3HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=0.8u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=1.12u l=0.12u
.ends XOR2M3HM
                                                           
.subckt XOR2M4HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.39u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
.ends XOR2M4HM
                                                           
.subckt XOR2M6HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.4u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=0.8u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.4u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.3u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=1.68u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.12u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.56u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.42u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=2.04u l=0.12u
.ends XOR2M6HM
                                                           
.subckt XOR2M8HM Z A B VDD VSS 
MN0 net01 A VSS VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN1 net02 B VSS VSS N_15_LL_EE2_UCFN w=1.12u l=0.12u
MN2 net03 net02 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN3 net03 A net04 VSS N_15_LL_EE2_UCFN w=0.52u l=0.12u
MN4 net02 net01 net04 VSS N_15_LL_EE2_UCFN w=0.48u l=0.12u
MN5 Z net04 VSS VSS N_15_LL_EE2_UCFN w=2.24u l=0.12u
MP0 VDD A net01 VDD P_15_LL_EE2_UCFN w=0.64u l=0.12u
MP1 VDD B net02 VDD P_15_LL_EE2_UCFN w=1.36u l=0.12u
MP2 VDD net02 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP3 net04 net01 net03 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP4 net04 A net02 VDD P_15_LL_EE2_UCFN w=0.72u l=0.12u
MP5 VDD net04 Z VDD P_15_LL_EE2_UCFN w=2.72u l=0.12u
.ends XOR2M8HM
                                                           
.subckt XOR3M0HM Z A B C VDD VSS 
MP17 VDD net126 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP23 VDD net153 net118 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP18 VDD net135 net94 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 net150 B net153 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP21 net94 net150 net126 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP22 net118 net141 net150 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP26 VDD C net135 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP27 net126 net138 net135 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP20 VDD A net153 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MP25 VDD net150 net138 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP24 VDD B net141 VDD P_15_LL_EE2_UCFN w=0.26u l=0.12u
MN17 Z net126 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN23 net147 net153 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN22 net150 B net147 VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN18 net129 net135 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN19 net153 net141 net150 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN21 net126 net138 net129 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN26 net135 C VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN24 net141 B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN27 net135 net150 net126 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net153 A VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN25 net138 net150 VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
.ends XOR3M0HM
                                                           
.subckt XOR3M1HM Z A B C VDD VSS 
MP17 VDD net126 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP23 VDD net153 net118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 VDD net135 net94 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 net150 B net153 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net94 net150 net126 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net118 net141 net150 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP26 VDD C net135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP27 net126 net138 net135 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP20 VDD A net153 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP25 VDD net150 net138 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP24 VDD B net141 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN17 Z net126 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN23 net147 net153 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN22 net150 B net147 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net129 net135 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN19 net153 net141 net150 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net126 net138 net129 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN26 net135 C VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN24 net141 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net135 net150 net126 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN20 net153 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN25 net138 net150 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends XOR3M1HM
                                                           
.subckt XOR3M2HM Z A B C VDD VSS 
MP17 VDD net126 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP23 VDD net153 net118 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP18 VDD net135 net94 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP19 net150 B net153 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP21 net94 net150 net126 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP22 net118 net141 net150 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP26 VDD C net135 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP27 net126 net138 net135 VDD P_15_LL_EE2_UCFN w=0.58u l=0.12u
MP20 VDD A net153 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP25 VDD net150 net138 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MP24 VDD B net141 VDD P_15_LL_EE2_UCFN w=0.35u l=0.12u
MN17 Z net126 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN23 net147 net153 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN22 net150 B net147 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN18 net129 net135 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN19 net153 net141 net150 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN21 net126 net138 net129 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN26 net135 C VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN24 net141 B VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN27 net135 net150 net126 VSS N_15_LL_EE2_UCFN w=0.46u l=0.12u
MN20 net153 A VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN25 net138 net150 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
.ends XOR3M2HM
                                                           
.subckt XOR3M4HM Z A B C VDD VSS 
MP17 VDD net126 Z VDD P_15_LL_EE2_UCFN w=1.28u l=0.12u
MP23 VDD net153 net118 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP18 VDD net135 net94 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP19 net150 B net153 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP21 net94 net150 net126 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP22 net118 net141 net150 VDD P_15_LL_EE2_UCFN w=0.34u l=0.12u
MP26 VDD C net135 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP27 net126 net138 net135 VDD P_15_LL_EE2_UCFN w=0.6u l=0.12u
MP20 VDD A net153 VDD P_15_LL_EE2_UCFN w=0.62u l=0.12u
MP25 VDD net150 net138 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP24 VDD B net141 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MN17 Z net126 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN23 net147 net153 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN22 net150 B net147 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN18 net129 net135 VSS VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN19 net153 net141 net150 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN21 net126 net138 net129 VSS N_15_LL_EE2_UCFN w=0.18u l=0.12u
MN26 net135 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN24 net141 B VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN27 net135 net150 net126 VSS N_15_LL_EE2_UCFN w=0.42u l=0.12u
MN20 net153 A VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN25 net138 net150 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
.ends XOR3M4HM
                                                           
.subckt XOR4M0HM Z A B C D VDD VSS 
MN14 Z net051 VSS VSS N_15_LL_EE2_UCFN w=0.31u l=0.12u
MN12 net083 net025 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN13 net080 net079 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN9 net0148 net080 net051 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net083 D net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0148 net081 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN8 net081 net079 net051 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net025 net022 net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net081 A net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 VSS net041 net014 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net081 net2 net041 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net022 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net025 C VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN1 net041 B VSS VSS N_15_LL_EE2_UCFN w=0.21u l=0.12u
MN0 net2 A VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MP14 VDD net051 Z VDD P_15_LL_EE2_UCFN w=0.38u l=0.12u
MP12 VDD net025 net083 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP11 net079 net022 net083 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 net079 D net025 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP13 VDD net079 net080 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net051 net080 net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 net051 net079 net0148 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD net081 net0148 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
MP6 net035 net2 net081 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP5 net035 net041 VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 net041 A net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD D net022 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD C net025 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP1 VDD B net041 VDD P_15_LL_EE2_UCFN w=0.29u l=0.12u
MP0 VDD A net2 VDD P_15_LL_EE2_UCFN w=0.25u l=0.12u
.ends XOR4M0HM
                                                           
.subckt XOR4M1HM Z A B C D VDD VSS 
MN14 Z net051 VSS VSS N_15_LL_EE2_UCFN w=0.39u l=0.12u
MN12 net083 net025 VSS VSS N_15_LL_EE2_UCFN w=0.24u l=0.12u
MN13 net080 net079 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN9 net0148 net080 net051 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN11 net083 D net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN7 net0148 net081 VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN8 net081 net079 net051 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN10 net025 net022 net079 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN6 net081 A net014 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN5 VSS net041 net014 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net081 net2 net041 VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN3 net022 D VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MN2 net025 C VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN1 net041 B VSS VSS N_15_LL_EE2_UCFN w=0.35u l=0.12u
MN0 net2 A VSS VSS N_15_LL_EE2_UCFN w=0.29u l=0.12u
MP14 VDD net051 Z VDD P_15_LL_EE2_UCFN w=0.48u l=0.12u
MP12 VDD net025 net083 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP11 net079 net022 net083 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP10 net079 D net025 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP13 VDD net079 net080 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net051 net080 net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 net051 net079 net0148 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD net081 net0148 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP6 net035 net2 net081 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP5 net035 net041 VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 net041 A net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP3 VDD D net022 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP2 VDD C net025 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP1 VDD B net041 VDD P_15_LL_EE2_UCFN w=0.49u l=0.12u
MP0 VDD A net2 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
.ends XOR4M1HM
                                                           
.subckt XOR4M2HM Z A B C D VDD VSS 
MN14 Z net051 VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN12 net083 net025 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN13 net080 net079 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN9 net0148 net080 net051 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN11 net083 D net079 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN7 net0148 net081 VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN8 net081 net079 net051 VSS N_15_LL_EE2_UCFN w=0.32u l=0.12u
MN10 net025 net022 net079 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN6 net081 A net014 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN5 VSS net041 net014 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net081 net2 net041 VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN3 net022 D VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MN2 net025 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN1 net041 B VSS VSS N_15_LL_EE2_UCFN w=0.56u l=0.12u
MN0 net2 A VSS VSS N_15_LL_EE2_UCFN w=0.37u l=0.12u
MP14 VDD net051 Z VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP12 VDD net025 net083 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP11 net079 net022 net083 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP10 net079 D net025 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP13 VDD net079 net080 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP8 net051 net080 net081 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 net051 net079 net0148 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP7 VDD net081 net0148 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP6 net035 net2 net081 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP5 net035 net041 VDD VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP4 net041 A net081 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP3 VDD D net022 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
MP2 VDD C net025 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP1 VDD B net041 VDD P_15_LL_EE2_UCFN w=0.68u l=0.12u
MP0 VDD A net2 VDD P_15_LL_EE2_UCFN w=0.46u l=0.12u
.ends XOR4M2HM
                                                           
.subckt XOR4M4HM Z A B C D VDD VSS 
MN14 Z net79 VSS VSS N_15_LL_EE2_UCFN w=1u l=0.12u
MN13 net10 D VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN12 net13 A VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN11 net16 C VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MN16 net0172 D net22 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN9 net22 net16 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN15 net0172 net10 net16 VSS N_15_LL_EE2_UCFN w=0.26u l=0.12u
MN7 net70 net0172 VSS VSS N_15_LL_EE2_UCFN w=0.19u l=0.12u
MN17 net79 net70 net37 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN18 net79 net0172 net47 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN4 net37 net47 VSS VSS N_15_LL_EE2_UCFN w=0.33u l=0.12u
MN3 net43 A net47 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN2 net43 net49 VSS VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN1 net49 net13 net47 VSS N_15_LL_EE2_UCFN w=0.28u l=0.12u
MN0 net49 B VSS VSS N_15_LL_EE2_UCFN w=0.5u l=0.12u
MP14 VDD net79 Z VDD P_15_LL_EE2_UCFN w=1.3u l=0.12u
MP13 VDD D net10 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP12 VDD A net13 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP11 VDD C net16 VDD P_15_LL_EE2_UCFN w=0.7u l=0.12u
MP16 net22 net10 net0172 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP9 VDD net16 net22 VDD P_15_LL_EE2_UCFN w=0.47u l=0.12u
MP15 net16 D net0172 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP7 VDD net0172 net70 VDD P_15_LL_EE2_UCFN w=0.28u l=0.12u
MP17 net37 net0172 net79 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP18 net47 net70 net79 VDD P_15_LL_EE2_UCFN w=0.33u l=0.12u
MP4 VDD net47 net37 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
MP3 net47 net13 net43 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP2 VDD net49 net43 VDD P_15_LL_EE2_UCFN w=0.32u l=0.12u
MP1 net47 A net49 VDD P_15_LL_EE2_UCFN w=0.36u l=0.12u
MP0 VDD B net49 VDD P_15_LL_EE2_UCFN w=0.65u l=0.12u
.ends XOR4M4HM
