module 接口列表阅读说明 #(
    parameter UDLY = 1
)(
endmodule