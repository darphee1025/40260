`timescale 1ns/1ps

`celldefine
module ADFM0HM( CO, S, A, B, CI , VDD, VSS);
inout VDD;
inout VSS;
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADFM0HM_func ADFM0HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));

   `else

	ADFM0HM_func ADFM0HM_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	ifnone
	// comb arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	ifnone
	// comb arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADFM1HM( CO, S, A, B, CI , VDD, VSS);
inout VDD;
inout VSS;
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADFM1HM_func ADFM1HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));

   `else

	ADFM1HM_func ADFM1HM_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	ifnone
	// comb arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	ifnone
	// comb arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADFM2HM( CO, S, A, B, CI , VDD, VSS);
inout VDD;
inout VSS;
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADFM2HM_func ADFM2HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));

   `else

	ADFM2HM_func ADFM2HM_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	ifnone
	// comb arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	ifnone
	// comb arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADFM4HM( CO, S, A, B, CI , VDD, VSS);
inout VDD;
inout VSS;
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADFM4HM_func ADFM4HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));

   `else

	ADFM4HM_func ADFM4HM_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	ifnone
	// comb arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	ifnone
	// comb arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADFM8HM( CO, S, A, B, CI , VDD, VSS);
inout VDD;
inout VSS;
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADFM8HM_func ADFM8HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));

   `else

	ADFM8HM_func ADFM8HM_inst(.CO(CO),.S(S),.A(A),.B(B),.CI(CI),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// comb arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// comb arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// comb arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	ifnone
	// comb arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	ifnone
	// comb arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc CI --> S
	 (CI => S) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADHM0HM( CO, S, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADHM0HM_func ADHM0HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ADHM0HM_func ADHM0HM_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADHM1HM( CO, S, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADHM1HM_func ADHM1HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ADHM1HM_func ADHM1HM_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADHM2HM( CO, S, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADHM2HM_func ADHM2HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ADHM2HM_func ADHM2HM_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADHM4HM( CO, S, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADHM4HM_func ADHM4HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ADHM4HM_func ADHM4HM_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADHM8HM( CO, S, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

	ADHM8HM_func ADHM8HM_behav_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ADHM8HM_func ADHM8HM_inst(.CO(CO),.S(S),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> CO
	 (A => CO) = (1.0,1.0);

	// comb arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M0HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M0HM_func AN2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M0HM_func AN2M0HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M12HM_func AN2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M12HM_func AN2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M16HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M16HM_func AN2M16HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M16HM_func AN2M16HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M1HM_func AN2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M1HM_func AN2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M2HM_func AN2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M2HM_func AN2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M4HM_func AN2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M4HM_func AN2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M6HM_func AN2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M6HM_func AN2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN2M8HM_func AN2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AN2M8HM_func AN2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M0HM_func AN3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M0HM_func AN3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M12HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M12HM_func AN3M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M12HM_func AN3M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M16HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M16HM_func AN3M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M16HM_func AN3M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M1HM_func AN3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M1HM_func AN3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M2HM_func AN3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M2HM_func AN3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M4HM_func AN3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M4HM_func AN3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M6HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M6HM_func AN3M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M6HM_func AN3M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN3M8HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN3M8HM_func AN3M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AN3M8HM_func AN3M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M0HM_func AN4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M0HM_func AN4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M12HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M12HM_func AN4M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M12HM_func AN4M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M16HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M16HM_func AN4M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M16HM_func AN4M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M1HM_func AN4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M1HM_func AN4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M2HM_func AN4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M2HM_func AN4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M4HM_func AN4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M4HM_func AN4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M6HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M6HM_func AN4M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M6HM_func AN4M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AN4M8HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AN4M8HM_func AN4M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	AN4M8HM_func AN4M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ANTHM( A );
input A;

endmodule
`endcelldefine

`celldefine
module AO211M0HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO211M0HM_func AO211M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO211M0HM_func AO211M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO211M1HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO211M1HM_func AO211M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO211M1HM_func AO211M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO211M2HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO211M2HM_func AO211M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO211M2HM_func AO211M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO211M4HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO211M4HM_func AO211M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO211M4HM_func AO211M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO211M8HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO211M8HM_func AO211M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO211M8HM_func AO211M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO21M0HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO21M0HM_func AO21M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO21M0HM_func AO21M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO21M1HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO21M1HM_func AO21M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO21M1HM_func AO21M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO21M2HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO21M2HM_func AO21M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO21M2HM_func AO21M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO21M4HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO21M4HM_func AO21M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO21M4HM_func AO21M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO21M8HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO21M8HM_func AO21M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO21M8HM_func AO21M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO221M0HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO221M0HM_func AO221M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO221M0HM_func AO221M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO221M1HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO221M1HM_func AO221M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO221M1HM_func AO221M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO221M2HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO221M2HM_func AO221M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO221M2HM_func AO221M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO221M4HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO221M4HM_func AO221M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO221M4HM_func AO221M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO221M8HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO221M8HM_func AO221M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AO221M8HM_func AO221M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO222M0HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO222M0HM_func AO222M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AO222M0HM_func AO222M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO222M1HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO222M1HM_func AO222M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AO222M1HM_func AO222M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO222M2HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO222M2HM_func AO222M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AO222M2HM_func AO222M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO222M4HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO222M4HM_func AO222M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AO222M4HM_func AO222M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO222M8HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO222M8HM_func AO222M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AO222M8HM_func AO222M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B10M0HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B10M0HM_func AO22B10M0HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B10M0HM_func AO22B10M0HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B10M1HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B10M1HM_func AO22B10M1HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B10M1HM_func AO22B10M1HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B10M2HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B10M2HM_func AO22B10M2HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B10M2HM_func AO22B10M2HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B10M4HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B10M4HM_func AO22B10M4HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B10M4HM_func AO22B10M4HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B10M8HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B10M8HM_func AO22B10M8HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B10M8HM_func AO22B10M8HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B11M0HM( Z, A1, B1, NA2, NB2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B11M0HM_func AO22B11M0HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B11M0HM_func AO22B11M0HM_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && NB2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B11M1HM( Z, A1, B1, NA2, NB2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B11M1HM_func AO22B11M1HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B11M1HM_func AO22B11M1HM_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && NB2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B11M2HM( Z, A1, B1, NA2, NB2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B11M2HM_func AO22B11M2HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B11M2HM_func AO22B11M2HM_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && NB2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B11M4HM( Z, A1, B1, NA2, NB2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B11M4HM_func AO22B11M4HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B11M4HM_func AO22B11M4HM_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && NB2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22B11M8HM( Z, A1, B1, NA2, NB2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22B11M8HM_func AO22B11M8HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));

   `else

	AO22B11M8HM_func AO22B11M8HM_inst(.Z(Z),.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && NB2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22M0HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22M0HM_func AO22M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO22M0HM_func AO22M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22M1HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22M1HM_func AO22M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO22M1HM_func AO22M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22M2HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22M2HM_func AO22M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO22M2HM_func AO22M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22M4HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22M4HM_func AO22M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO22M4HM_func AO22M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO22M8HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO22M8HM_func AO22M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO22M8HM_func AO22M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO31M0HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO31M0HM_func AO31M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO31M0HM_func AO31M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO31M1HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO31M1HM_func AO31M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO31M1HM_func AO31M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO31M2HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO31M2HM_func AO31M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO31M2HM_func AO31M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO31M4HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO31M4HM_func AO31M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO31M4HM_func AO31M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO31M8HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO31M8HM_func AO31M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AO31M8HM_func AO31M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO32M0HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO32M0HM_func AO32M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO32M0HM_func AO32M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO32M1HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO32M1HM_func AO32M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO32M1HM_func AO32M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO32M2HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO32M2HM_func AO32M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO32M2HM_func AO32M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO32M4HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO32M4HM_func AO32M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO32M4HM_func AO32M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO32M8HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO32M8HM_func AO32M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AO32M8HM_func AO32M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO33M0HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO33M0HM_func AO33M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AO33M0HM_func AO33M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO33M1HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO33M1HM_func AO33M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AO33M1HM_func AO33M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO33M2HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO33M2HM_func AO33M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AO33M2HM_func AO33M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO33M4HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO33M4HM_func AO33M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AO33M4HM_func AO33M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AO33M8HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AO33M8HM_func AO33M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AO33M8HM_func AO33M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI211M0HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI211M0HM_func AOI211M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI211M0HM_func AOI211M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI211M1HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI211M1HM_func AOI211M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI211M1HM_func AOI211M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI211M2HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI211M2HM_func AOI211M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI211M2HM_func AOI211M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI211M4HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI211M4HM_func AOI211M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI211M4HM_func AOI211M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI211M8HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI211M8HM_func AOI211M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI211M8HM_func AOI211M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B01M0HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M0HM_func AOI21B01M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B01M0HM_func AOI21B01M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B01M1HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M1HM_func AOI21B01M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B01M1HM_func AOI21B01M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B01M2HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M2HM_func AOI21B01M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B01M2HM_func AOI21B01M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B01M4HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M4HM_func AOI21B01M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B01M4HM_func AOI21B01M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B01M8HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M8HM_func AOI21B01M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B01M8HM_func AOI21B01M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B10M0HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M0HM_func AOI21B10M0HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B10M0HM_func AOI21B10M0HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B10M1HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M1HM_func AOI21B10M1HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B10M1HM_func AOI21B10M1HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B10M2HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M2HM_func AOI21B10M2HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B10M2HM_func AOI21B10M2HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B10M4HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M4HM_func AOI21B10M4HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B10M4HM_func AOI21B10M4HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B10M8HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M8HM_func AOI21B10M8HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B10M8HM_func AOI21B10M8HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B20M0HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M0HM_func AOI21B20M0HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B20M0HM_func AOI21B20M0HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B20M1HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M1HM_func AOI21B20M1HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B20M1HM_func AOI21B20M1HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B20M2HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M2HM_func AOI21B20M2HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B20M2HM_func AOI21B20M2HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B20M4HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M4HM_func AOI21B20M4HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B20M4HM_func AOI21B20M4HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21B20M8HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M8HM_func AOI21B20M8HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI21B20M8HM_func AOI21B20M8HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M0HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M0HM_func AOI21M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M0HM_func AOI21M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M1HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M1HM_func AOI21M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M1HM_func AOI21M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M2HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M2HM_func AOI21M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M2HM_func AOI21M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M3HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M3HM_func AOI21M3HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M3HM_func AOI21M3HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M4HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M4HM_func AOI21M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M4HM_func AOI21M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M6HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M6HM_func AOI21M6HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M6HM_func AOI21M6HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI21M8HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI21M8HM_func AOI21M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI21M8HM_func AOI21M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI221M0HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI221M0HM_func AOI221M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI221M0HM_func AOI221M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI221M1HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI221M1HM_func AOI221M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI221M1HM_func AOI221M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI221M2HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI221M2HM_func AOI221M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI221M2HM_func AOI221M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI221M4HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI221M4HM_func AOI221M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI221M4HM_func AOI221M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI221M8HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI221M8HM_func AOI221M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	AOI221M8HM_func AOI221M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI222M0HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI222M0HM_func AOI222M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AOI222M0HM_func AOI222M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI222M1HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI222M1HM_func AOI222M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AOI222M1HM_func AOI222M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI222M2HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI222M2HM_func AOI222M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AOI222M2HM_func AOI222M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI222M4HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI222M4HM_func AOI222M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AOI222M4HM_func AOI222M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI222M8HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI222M8HM_func AOI222M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	AOI222M8HM_func AOI222M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22B20M0HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M0HM_func AOI22B20M0HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22B20M0HM_func AOI22B20M0HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22B20M1HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M1HM_func AOI22B20M1HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22B20M1HM_func AOI22B20M1HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22B20M2HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M2HM_func AOI22B20M2HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22B20M2HM_func AOI22B20M2HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22B20M4HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M4HM_func AOI22B20M4HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22B20M4HM_func AOI22B20M4HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22B20M8HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M8HM_func AOI22B20M8HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22B20M8HM_func AOI22B20M8HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22M0HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22M0HM_func AOI22M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22M0HM_func AOI22M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22M1HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22M1HM_func AOI22M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22M1HM_func AOI22M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22M2HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22M2HM_func AOI22M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22M2HM_func AOI22M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22M4HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22M4HM_func AOI22M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22M4HM_func AOI22M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI22M8HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI22M8HM_func AOI22M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI22M8HM_func AOI22M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI31M0HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI31M0HM_func AOI31M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI31M0HM_func AOI31M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI31M1HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI31M1HM_func AOI31M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI31M1HM_func AOI31M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI31M2HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI31M2HM_func AOI31M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI31M2HM_func AOI31M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI31M4HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI31M4HM_func AOI31M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI31M4HM_func AOI31M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI31M8HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI31M8HM_func AOI31M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	AOI31M8HM_func AOI31M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI32M0HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI32M0HM_func AOI32M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI32M0HM_func AOI32M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI32M1HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI32M1HM_func AOI32M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI32M1HM_func AOI32M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI32M2HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI32M2HM_func AOI32M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI32M2HM_func AOI32M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI32M4HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI32M4HM_func AOI32M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI32M4HM_func AOI32M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI32M8HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI32M8HM_func AOI32M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	AOI32M8HM_func AOI32M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI33M0HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI33M0HM_func AOI33M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AOI33M0HM_func AOI33M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI33M1HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI33M1HM_func AOI33M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AOI33M1HM_func AOI33M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI33M2HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI33M2HM_func AOI33M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AOI33M2HM_func AOI33M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI33M4HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI33M4HM_func AOI33M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AOI33M4HM_func AOI33M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module AOI33M8HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	AOI33M8HM_func AOI33M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	AOI33M8HM_func AOI33M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BHDM1HM( Z, VDD, VSS);
inout VDD;
inout VSS;
inout Z;

    // Busholder.
wire io_wire, Z_org;

bufif1 (Z_org, 1'bx, (VDD != 1'b1 || VSS != 1'b0 ));
bufif0 (Z_org, Z, (VDD != 1'b1 || VSS != 1'b0 ));
  buf(weak0,weak1) SMC_I0(Z, io_wire);
  buf              SMC_I1(io_wire, Z_org);
 
endmodule
`endcelldefine

`celldefine
module BUFM10HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM10HM_func BUFM10HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM10HM_func BUFM10HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM12HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM12HM_func BUFM12HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM12HM_func BUFM12HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM14HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM14HM_func BUFM14HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM14HM_func BUFM14HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM16HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM16HM_func BUFM16HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM16HM_func BUFM16HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM18HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM18HM_func BUFM18HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM18HM_func BUFM18HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM20HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM20HM_func BUFM20HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM20HM_func BUFM20HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM24HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM24HM_func BUFM24HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM24HM_func BUFM24HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM28HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM28HM_func BUFM28HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM28HM_func BUFM28HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM2HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM2HM_func BUFM2HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM2HM_func BUFM2HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM32HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM32HM_func BUFM32HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM32HM_func BUFM32HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM36HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM36HM_func BUFM36HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM36HM_func BUFM36HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM3HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM3HM_func BUFM3HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM3HM_func BUFM3HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM40HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM40HM_func BUFM40HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM40HM_func BUFM40HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM48HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM48HM_func BUFM48HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM48HM_func BUFM48HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM4HM_func BUFM4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM4HM_func BUFM4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM5HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM5HM_func BUFM5HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM5HM_func BUFM5HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM6HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM6HM_func BUFM6HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM6HM_func BUFM6HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFM8HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFM8HM_func BUFM8HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	BUFM8HM_func BUFM8HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM12HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM12HM_func BUFTM12HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM12HM_func BUFTM12HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM16HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM16HM_func BUFTM16HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM16HM_func BUFTM16HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM1HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM1HM_func BUFTM1HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM1HM_func BUFTM1HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM20HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM20HM_func BUFTM20HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM20HM_func BUFTM20HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM24HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM24HM_func BUFTM24HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM24HM_func BUFTM24HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM2HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM2HM_func BUFTM2HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM2HM_func BUFTM2HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM3HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM3HM_func BUFTM3HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM3HM_func BUFTM3HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM4HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM4HM_func BUFTM4HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM4HM_func BUFTM4HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM6HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM6HM_func BUFTM6HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM6HM_func BUFTM6HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module BUFTM8HM( Z, A, E , VDD, VSS);
inout VDD;
inout VSS;
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	BUFTM8HM_func BUFTM8HM_behav_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));

   `else

	BUFTM8HM_func BUFTM8HM_inst(.Z(Z),.A(A),.E(E),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M12HM_func CKAN2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M12HM_func CKAN2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M16HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M16HM_func CKAN2M16HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M16HM_func CKAN2M16HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M2HM_func CKAN2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M2HM_func CKAN2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M3HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M3HM_func CKAN2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M3HM_func CKAN2M3HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M4HM_func CKAN2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M4HM_func CKAN2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M6HM_func CKAN2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M6HM_func CKAN2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKAN2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKAN2M8HM_func CKAN2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKAN2M8HM_func CKAN2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM12HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM12HM_func CKBUFM12HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM12HM_func CKBUFM12HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM16HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM16HM_func CKBUFM16HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM16HM_func CKBUFM16HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM1HM_func CKBUFM1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM1HM_func CKBUFM1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM20HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM20HM_func CKBUFM20HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM20HM_func CKBUFM20HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM24HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM24HM_func CKBUFM24HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM24HM_func CKBUFM24HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM2HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM2HM_func CKBUFM2HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM2HM_func CKBUFM2HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM32HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM32HM_func CKBUFM32HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM32HM_func CKBUFM32HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM3HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM3HM_func CKBUFM3HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM3HM_func CKBUFM3HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM40HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM40HM_func CKBUFM40HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM40HM_func CKBUFM40HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM48HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM48HM_func CKBUFM48HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM48HM_func CKBUFM48HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM4HM_func CKBUFM4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM4HM_func CKBUFM4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM6HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM6HM_func CKBUFM6HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM6HM_func CKBUFM6HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKBUFM8HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKBUFM8HM_func CKBUFM8HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKBUFM8HM_func CKBUFM8HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM12HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM12HM_func CKINVM12HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM12HM_func CKINVM12HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM16HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM16HM_func CKINVM16HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM16HM_func CKINVM16HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM1HM_func CKINVM1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM1HM_func CKINVM1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM20HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM20HM_func CKINVM20HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM20HM_func CKINVM20HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM24HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM24HM_func CKINVM24HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM24HM_func CKINVM24HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM2HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM2HM_func CKINVM2HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM2HM_func CKINVM2HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM32HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM32HM_func CKINVM32HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM32HM_func CKINVM32HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM3HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM3HM_func CKINVM3HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM3HM_func CKINVM3HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM40HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM40HM_func CKINVM40HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM40HM_func CKINVM40HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM48HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM48HM_func CKINVM48HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM48HM_func CKINVM48HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM4HM_func CKINVM4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM4HM_func CKINVM4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM6HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM6HM_func CKINVM6HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM6HM_func CKINVM6HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKINVM8HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKINVM8HM_func CKINVM8HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	CKINVM8HM_func CKINVM8HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKMUX2M12HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M12HM_func CKMUX2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	CKMUX2M12HM_func CKMUX2M12HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKMUX2M2HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M2HM_func CKMUX2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	CKMUX2M2HM_func CKMUX2M2HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKMUX2M3HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M3HM_func CKMUX2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	CKMUX2M3HM_func CKMUX2M3HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKMUX2M4HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M4HM_func CKMUX2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	CKMUX2M4HM_func CKMUX2M4HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKMUX2M6HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M6HM_func CKMUX2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	CKMUX2M6HM_func CKMUX2M6HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKMUX2M8HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M8HM_func CKMUX2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	CKMUX2M8HM_func CKMUX2M8HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKND2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKND2M12HM_func CKND2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKND2M12HM_func CKND2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKND2M16HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKND2M16HM_func CKND2M16HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKND2M16HM_func CKND2M16HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKND2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKND2M2HM_func CKND2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKND2M2HM_func CKND2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKND2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKND2M4HM_func CKND2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKND2M4HM_func CKND2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKND2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKND2M6HM_func CKND2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKND2M6HM_func CKND2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKND2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKND2M8HM_func CKND2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKND2M8HM_func CKND2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKXOR2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M12HM_func CKXOR2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKXOR2M12HM_func CKXOR2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKXOR2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M1HM_func CKXOR2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKXOR2M1HM_func CKXOR2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKXOR2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M2HM_func CKXOR2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKXOR2M2HM_func CKXOR2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKXOR2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M4HM_func CKXOR2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKXOR2M4HM_func CKXOR2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module CKXOR2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M8HM_func CKXOR2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	CKXOR2M8HM_func CKXOR2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL1M1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL1M1HM_func DEL1M1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL1M1HM_func DEL1M1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL1M4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL1M4HM_func DEL1M4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL1M4HM_func DEL1M4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL2M1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL2M1HM_func DEL2M1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL2M1HM_func DEL2M1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL2M4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL2M4HM_func DEL2M4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL2M4HM_func DEL2M4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL3M1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL3M1HM_func DEL3M1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL3M1HM_func DEL3M1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL3M4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL3M4HM_func DEL3M4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL3M4HM_func DEL3M4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL4M1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL4M1HM_func DEL4M1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL4M1HM_func DEL4M1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DEL4M4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	DEL4M4HM_func DEL4M4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	DEL4M4HM_func DEL4M4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCM1HM( Q, QB, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCM1HM_func DFCM1HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCM1HM_func DFCM1HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCM2HM( Q, QB, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCM2HM_func DFCM2HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCM2HM_func DFCM2HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCM4HM( Q, QB, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCM4HM_func DFCM4HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCM4HM_func DFCM4HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCM8HM( Q, QB, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCM8HM_func DFCM8HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCM8HM_func DFCM8HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQM1HM( Q, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQM1HM_func DFCQM1HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCQM1HM_func DFCQM1HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQM2HM( Q, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQM2HM_func DFCQM2HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCQM2HM_func DFCQM2HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQM4HM( Q, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQM4HM_func DFCQM4HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCQM4HM_func DFCQM4HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQM8HM( Q, CKB, D , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQM8HM_func DFCQM8HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	DFCQM8HM_func DFCQM8HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQRSM1HM( Q, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM1HM_func DFCQRSM1HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCQRSM1HM_func DFCQRSM1HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQRSM2HM( Q, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM2HM_func DFCQRSM2HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCQRSM2HM_func DFCQRSM2HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQRSM4HM( Q, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM4HM_func DFCQRSM4HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCQRSM4HM_func DFCQRSM4HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCQRSM8HM( Q, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM8HM_func DFCQRSM8HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCQRSM8HM_func DFCQRSM8HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCRSM1HM( Q, QB, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCRSM1HM_func DFCRSM1HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCRSM1HM_func DFCRSM1HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCRSM2HM( Q, QB, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCRSM2HM_func DFCRSM2HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCRSM2HM_func DFCRSM2HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCRSM4HM( Q, QB, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCRSM4HM_func DFCRSM4HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCRSM4HM_func DFCRSM4HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFCRSM8HM( Q, QB, CKB, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFCRSM8HM_func DFCRSM8HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFCRSM8HM_func DFCRSM8HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CKB$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CKB$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CKB_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CKB$delay);


	and MGM_G16(ENABLE_CKB_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CKB$delay);


	and MGM_G18(ENABLE_CKB_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CKB$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CKB_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CKB$delay);


	and MGM_G23(ENABLE_NOT_CKB_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CKB_AND_NOT_D,MGM_W14,CKB$delay);


	and MGM_G26(ENABLE_CKB_AND_D,D$delay,CKB$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CKB$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CKB$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CKB_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CKB$delay);


	and MGM_G37(ENABLE_CKB_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CKB$delay);


	and MGM_G39(ENABLE_CKB_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEM1HM( Q, QB, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEM1HM_func DFEM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEM1HM_func DFEM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEM2HM( Q, QB, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEM2HM_func DFEM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEM2HM_func DFEM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEM4HM( Q, QB, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEM4HM_func DFEM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEM4HM_func DFEM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEM8HM( Q, QB, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEM8HM_func DFEM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEM8HM_func DFEM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQM1HM( Q, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQM1HM_func DFEQM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEQM1HM_func DFEQM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQM2HM( Q, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQM2HM_func DFEQM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEQM2HM_func DFEQM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQM4HM( Q, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQM4HM_func DFEQM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEQM4HM_func DFEQM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQM8HM( Q, CK, D, E , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQM8HM_func DFEQM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	DFEQM8HM_func DFEQM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_E,E$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_E,E$delay,D$delay);


	buf MGM_G3(ENABLE_E,E$delay);


	not MGM_G4(ENABLE_NOT_D,D$delay);


	buf MGM_G5(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		posedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1),
		negedge E &&& (ENABLE_NOT_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		posedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D === 1'b1),
		negedge E &&& (ENABLE_D === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQRM1HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQRM1HM_func DFEQRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQRM1HM_func DFEQRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQRM2HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQRM2HM_func DFEQRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQRM2HM_func DFEQRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQRM4HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQRM4HM_func DFEQRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQRM4HM_func DFEQRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQRM8HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQRM8HM_func DFEQRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQRM8HM_func DFEQRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQZRM1HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM1HM_func DFEQZRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQZRM1HM_func DFEQZRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQZRM2HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM2HM_func DFEQZRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQZRM2HM_func DFEQZRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQZRM4HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM4HM_func DFEQZRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQZRM4HM_func DFEQZRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEQZRM8HM( Q, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM8HM_func DFEQZRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEQZRM8HM_func DFEQZRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFERM1HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFERM1HM_func DFERM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFERM1HM_func DFERM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFERM2HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFERM2HM_func DFERM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFERM2HM_func DFERM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFERM4HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFERM4HM_func DFERM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFERM4HM_func DFERM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFERM8HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFERM8HM_func DFERM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFERM8HM_func DFERM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,E$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W1);


	and MGM_G3(MGM_W2,E$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W2);


	and MGM_G5(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G6(MGM_W3,D$delay);


	and MGM_G7(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W3);


	and MGM_G8(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G9(ENABLE_E,E$delay);


	not MGM_G10(MGM_W4,CK$delay);


	not MGM_G11(MGM_W5,D$delay);


	and MGM_G12(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G13(MGM_W7,E$delay);


	and MGM_G14(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E,MGM_W7,MGM_W6);


	not MGM_G15(MGM_W8,CK$delay);


	not MGM_G16(MGM_W9,D$delay);


	and MGM_G17(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G18(ENABLE_NOT_CK_AND_NOT_D_AND_E,E$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	and MGM_G20(MGM_W12,D$delay,MGM_W11);


	not MGM_G21(MGM_W13,E$delay);


	and MGM_G22(ENABLE_NOT_CK_AND_D_AND_NOT_E,MGM_W13,MGM_W12);


	not MGM_G23(MGM_W14,CK$delay);


	and MGM_G24(MGM_W15,D$delay,MGM_W14);


	and MGM_G25(ENABLE_NOT_CK_AND_D_AND_E,E$delay,MGM_W15);


	not MGM_G26(MGM_W16,D$delay);


	and MGM_G27(MGM_W17,MGM_W16,CK$delay);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_CK_AND_NOT_D_AND_NOT_E,MGM_W18,MGM_W17);


	not MGM_G30(MGM_W19,D$delay);


	and MGM_G31(MGM_W20,MGM_W19,CK$delay);


	and MGM_G32(ENABLE_CK_AND_NOT_D_AND_E,E$delay,MGM_W20);


	and MGM_G33(MGM_W21,D$delay,CK$delay);


	not MGM_G34(MGM_W22,E$delay);


	and MGM_G35(ENABLE_CK_AND_D_AND_NOT_E,MGM_W22,MGM_W21);


	and MGM_G36(MGM_W23,D$delay,CK$delay);


	and MGM_G37(ENABLE_CK_AND_D_AND_E,E$delay,MGM_W23);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_E === 1'b1),
		posedge CK &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEZRM1HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEZRM1HM_func DFEZRM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEZRM1HM_func DFEZRM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEZRM2HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEZRM2HM_func DFEZRM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEZRM2HM_func DFEZRM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEZRM4HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEZRM4HM_func DFEZRM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEZRM4HM_func DFEZRM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFEZRM8HM( Q, QB, CK, D, E, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFEZRM8HM_func DFEZRM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	DFEZRM8HM_func DFEZRM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	and MGM_G6(MGM_W5,E$delay,MGM_W4);


	not MGM_G7(MGM_W6,RB$delay);


	and MGM_G8(ENABLE_NOT_D_AND_E_AND_NOT_RB,MGM_W6,MGM_W5);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,E$delay,MGM_W7);


	and MGM_G11(ENABLE_NOT_D_AND_E_AND_RB,RB$delay,MGM_W8);


	not MGM_G12(MGM_W9,E$delay);


	and MGM_G13(MGM_W10,MGM_W9,D$delay);


	not MGM_G14(MGM_W11,RB$delay);


	and MGM_G15(ENABLE_D_AND_NOT_E_AND_NOT_RB,MGM_W11,MGM_W10);


	and MGM_G16(MGM_W12,E$delay,D$delay);


	not MGM_G17(MGM_W13,RB$delay);


	and MGM_G18(ENABLE_D_AND_E_AND_NOT_RB,MGM_W13,MGM_W12);


	and MGM_G19(MGM_W14,E$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_E_AND_RB,RB$delay,MGM_W14);


	and MGM_G21(ENABLE_E_AND_RB,RB$delay,E$delay);


	not MGM_G22(MGM_W15,D$delay);


	and MGM_G23(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W15);


	and MGM_G24(ENABLE_D_AND_RB,RB$delay,D$delay);


	not MGM_G25(MGM_W16,D$delay);


	not MGM_G26(MGM_W17,E$delay);


	and MGM_G27(ENABLE_NOT_D_AND_NOT_E,MGM_W17,MGM_W16);


	not MGM_G28(MGM_W18,E$delay);


	and MGM_G29(ENABLE_D_AND_NOT_E,MGM_W18,D$delay);


	and MGM_G30(ENABLE_D_AND_E,E$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFM1HM( Q, QB, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFM1HM_func DFM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFM1HM_func DFM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFM2HM( Q, QB, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFM2HM_func DFM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFM2HM_func DFM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFM4HM( Q, QB, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFM4HM_func DFM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFM4HM_func DFM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFM8HM( Q, QB, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFM8HM_func DFM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFM8HM_func DFM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMM1HM( Q, QB, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMM1HM_func DFMM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMM1HM_func DFMM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMM2HM( Q, QB, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMM2HM_func DFMM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMM2HM_func DFMM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMM4HM( Q, QB, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMM4HM_func DFMM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMM4HM_func DFMM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMM8HM( Q, QB, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMM8HM_func DFMM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMM8HM_func DFMM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMQM1HM( Q, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMQM1HM_func DFMQM1HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMQM1HM_func DFMQM1HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMQM2HM( Q, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMQM2HM_func DFMQM2HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMQM2HM_func DFMQM2HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMQM4HM( Q, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMQM4HM_func DFMQM4HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMQM4HM_func DFMQM4HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFMQM8HM( Q, CK, D1, D2, S , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFMQM8HM_func DFMQM8HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	DFMQM8HM_func DFMQM8HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D1$delay);


	not MGM_G6(MGM_W5,D2$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_S,S$delay,MGM_W6);


	not MGM_G9(MGM_W7,D1$delay);


	and MGM_G10(MGM_W8,D2$delay,MGM_W7);


	not MGM_G11(MGM_W9,S$delay);


	and MGM_G12(ENABLE_NOT_D1_AND_D2_AND_NOT_S,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D1$delay);


	and MGM_G14(MGM_W11,D2$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D1_AND_D2_AND_S,S$delay,MGM_W11);


	not MGM_G16(MGM_W12,D2$delay);


	and MGM_G17(MGM_W13,MGM_W12,D1$delay);


	not MGM_G18(MGM_W14,S$delay);


	and MGM_G19(ENABLE_D1_AND_NOT_D2_AND_NOT_S,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,D2$delay);


	and MGM_G21(MGM_W16,MGM_W15,D1$delay);


	and MGM_G22(ENABLE_D1_AND_NOT_D2_AND_S,S$delay,MGM_W16);


	and MGM_G23(MGM_W17,D2$delay,D1$delay);


	not MGM_G24(MGM_W18,S$delay);


	and MGM_G25(ENABLE_D1_AND_D2_AND_NOT_S,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,D2$delay,D1$delay);


	and MGM_G27(ENABLE_D1_AND_D2_AND_S,S$delay,MGM_W19);


	not MGM_G28(MGM_W20,D2$delay);


	and MGM_G29(ENABLE_NOT_D2_AND_S,S$delay,MGM_W20);


	and MGM_G30(ENABLE_D2_AND_S,S$delay,D2$delay);


	not MGM_G31(MGM_W21,D1$delay);


	not MGM_G32(MGM_W22,S$delay);


	and MGM_G33(ENABLE_NOT_D1_AND_NOT_S,MGM_W22,MGM_W21);


	not MGM_G34(MGM_W23,S$delay);


	and MGM_G35(ENABLE_D1_AND_NOT_S,MGM_W23,D1$delay);


	not MGM_G36(MGM_W24,D1$delay);


	and MGM_G37(ENABLE_NOT_D1_AND_D2,D2$delay,MGM_W24);


	not MGM_G38(MGM_W25,D2$delay);


	and MGM_G39(ENABLE_D1_AND_NOT_D2,MGM_W25,D1$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2 === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQM1HM( Q, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQM1HM_func DFQM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFQM1HM_func DFQM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQM2HM( Q, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQM2HM_func DFQM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFQM2HM_func DFQM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQM4HM( Q, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQM4HM_func DFQM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFQM4HM_func DFQM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQM8HM( Q, CK, D , VDD, VSS);
inout VDD;
inout VSS;
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQM8HM_func DFQM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	DFQM8HM_func DFQM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRM1HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRM1HM_func DFQRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQRM1HM_func DFQRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRM2HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRM2HM_func DFQRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQRM2HM_func DFQRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRM4HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRM4HM_func DFQRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQRM4HM_func DFQRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRM8HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRM8HM_func DFQRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQRM8HM_func DFQRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRSM1HM( Q, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRSM1HM_func DFQRSM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFQRSM1HM_func DFQRSM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRSM2HM( Q, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRSM2HM_func DFQRSM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFQRSM2HM_func DFQRSM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRSM4HM( Q, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRSM4HM_func DFQRSM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFQRSM4HM_func DFQRSM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQRSM8HM( Q, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQRSM8HM_func DFQRSM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFQRSM8HM_func DFQRSM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQSM1HM( Q, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQSM1HM_func DFQSM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFQSM1HM_func DFQSM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQSM2HM( Q, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQSM2HM_func DFQSM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFQSM2HM_func DFQSM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQSM4HM( Q, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQSM4HM_func DFQSM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFQSM4HM_func DFQSM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQSM8HM( Q, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQSM8HM_func DFQSM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFQSM8HM_func DFQSM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQZRM1HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQZRM1HM_func DFQZRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQZRM1HM_func DFQZRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQZRM2HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQZRM2HM_func DFQZRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQZRM2HM_func DFQZRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQZRM4HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQZRM4HM_func DFQZRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQZRM4HM_func DFQZRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFQZRM8HM( Q, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFQZRM8HM_func DFQZRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFQZRM8HM_func DFQZRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRM1HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRM1HM_func DFRM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFRM1HM_func DFRM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRM2HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRM2HM_func DFRM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFRM2HM_func DFRM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRM4HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRM4HM_func DFRM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFRM4HM_func DFRM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRM8HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRM8HM_func DFRM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFRM8HM_func DFRM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_RB,RB$delay,D$delay);


	buf MGM_G3(ENABLE_RB,RB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRSM1HM( Q, QB, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRSM1HM_func DFRSM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFRSM1HM_func DFRSM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRSM2HM( Q, QB, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRSM2HM_func DFRSM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFRSM2HM_func DFRSM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRSM4HM( Q, QB, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRSM4HM_func DFRSM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFRSM4HM_func DFRSM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFRSM8HM( Q, QB, CK, D, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFRSM8HM_func DFRSM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	DFRSM8HM_func DFRSM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G3(MGM_W2,RB$delay,D$delay);


	and MGM_G4(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	and MGM_G5(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,CK$delay);


	not MGM_G8(MGM_W4,D$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,CK$delay);


	and MGM_G12(MGM_W7,D$delay,MGM_W6);


	and MGM_G13(ENABLE_NOT_CK_AND_D_AND_SB,SB$delay,MGM_W7);


	not MGM_G14(MGM_W8,D$delay);


	and MGM_G15(MGM_W9,MGM_W8,CK$delay);


	and MGM_G16(ENABLE_CK_AND_NOT_D_AND_SB,SB$delay,MGM_W9);


	and MGM_G17(MGM_W10,D$delay,CK$delay);


	and MGM_G18(ENABLE_CK_AND_D_AND_SB,SB$delay,MGM_W10);


	not MGM_G19(MGM_W11,CK$delay);


	not MGM_G20(MGM_W12,D$delay);


	and MGM_G21(ENABLE_NOT_CK_AND_NOT_D,MGM_W12,MGM_W11);


	not MGM_G22(MGM_W13,CK$delay);


	and MGM_G23(ENABLE_NOT_CK_AND_D,D$delay,MGM_W13);


	not MGM_G24(MGM_W14,D$delay);


	and MGM_G25(ENABLE_CK_AND_NOT_D,MGM_W14,CK$delay);


	and MGM_G26(ENABLE_CK_AND_D,D$delay,CK$delay);


	buf MGM_G27(ENABLE_RB,RB$delay);


	not MGM_G28(MGM_W15,CK$delay);


	not MGM_G29(MGM_W16,D$delay);


	and MGM_G30(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G31(ENABLE_NOT_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W17);


	not MGM_G32(MGM_W18,CK$delay);


	and MGM_G33(MGM_W19,D$delay,MGM_W18);


	and MGM_G34(ENABLE_NOT_CK_AND_D_AND_RB,RB$delay,MGM_W19);


	not MGM_G35(MGM_W20,D$delay);


	and MGM_G36(MGM_W21,MGM_W20,CK$delay);


	and MGM_G37(ENABLE_CK_AND_NOT_D_AND_RB,RB$delay,MGM_W21);


	and MGM_G38(MGM_W22,D$delay,CK$delay);


	and MGM_G39(ENABLE_CK_AND_D_AND_RB,RB$delay,MGM_W22);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFSM1HM( Q, QB, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFSM1HM_func DFSM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFSM1HM_func DFSM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFSM2HM( Q, QB, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFSM2HM_func DFSM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFSM2HM_func DFSM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFSM4HM( Q, QB, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFSM4HM_func DFSM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFSM4HM_func DFSM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFSM8HM( Q, QB, CK, D, SB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFSM8HM_func DFSM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	DFSM8HM_func DFSM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(ENABLE_NOT_D_AND_SB,SB$delay,MGM_W0);


	and MGM_G2(ENABLE_D_AND_SB,SB$delay,D$delay);


	buf MGM_G3(ENABLE_SB,SB$delay);


	not MGM_G4(MGM_W1,CK$delay);


	not MGM_G5(MGM_W2,D$delay);


	and MGM_G6(ENABLE_NOT_CK_AND_NOT_D,MGM_W2,MGM_W1);


	not MGM_G7(MGM_W3,CK$delay);


	and MGM_G8(ENABLE_NOT_CK_AND_D,D$delay,MGM_W3);


	not MGM_G9(MGM_W4,D$delay);


	and MGM_G10(ENABLE_CK_AND_NOT_D,MGM_W4,CK$delay);


	and MGM_G11(ENABLE_CK_AND_D,D$delay,CK$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D === 1'b1)
		,1.0,0,notifier);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFZRM1HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFZRM1HM_func DFZRM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFZRM1HM_func DFZRM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFZRM2HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFZRM2HM_func DFZRM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFZRM2HM_func DFZRM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFZRM4HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFZRM4HM_func DFZRM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFZRM4HM_func DFZRM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module DFZRM8HM( Q, QB, CK, D, RB , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	DFZRM8HM_func DFZRM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	DFZRM8HM_func DFZRM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(ENABLE_NOT_D_AND_NOT_RB,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,D$delay);


	and MGM_G4(ENABLE_NOT_D_AND_RB,RB$delay,MGM_W2);


	not MGM_G5(MGM_W3,RB$delay);


	and MGM_G6(ENABLE_D_AND_NOT_RB,MGM_W3,D$delay);


	and MGM_G7(ENABLE_D_AND_RB,RB$delay,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM0HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM0HM_func INVM0HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM0HM_func INVM0HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM10HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM10HM_func INVM10HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM10HM_func INVM10HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM12HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM12HM_func INVM12HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM12HM_func INVM12HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM14HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM14HM_func INVM14HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM14HM_func INVM14HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM16HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM16HM_func INVM16HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM16HM_func INVM16HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM18HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM18HM_func INVM18HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM18HM_func INVM18HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM1HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM1HM_func INVM1HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM1HM_func INVM1HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM20HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM20HM_func INVM20HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM20HM_func INVM20HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM24HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM24HM_func INVM24HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM24HM_func INVM24HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM28HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM28HM_func INVM28HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM28HM_func INVM28HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM2HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM2HM_func INVM2HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM2HM_func INVM2HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM32HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM32HM_func INVM32HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM32HM_func INVM32HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM36HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM36HM_func INVM36HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM36HM_func INVM36HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM3HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM3HM_func INVM3HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM3HM_func INVM3HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM40HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM40HM_func INVM40HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM40HM_func INVM40HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM48HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM48HM_func INVM48HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM48HM_func INVM48HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM4HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM4HM_func INVM4HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM4HM_func INVM4HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM5HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM5HM_func INVM5HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM5HM_func INVM5HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM6HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM6HM_func INVM6HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM6HM_func INVM6HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module INVM8HM( Z, A , VDD, VSS);
inout VDD;
inout VSS;
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	INVM8HM_func INVM8HM_behav_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));

   `else

	INVM8HM_func INVM8HM_inst(.Z(Z),.A(A),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACM0HM( Q, QB, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACM0HM_func LACM0HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	LACM0HM_func LACM0HM_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D);


	buf MGM_G1(ENABLE_D,D);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 


   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACM1HM( Q, QB, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACM1HM_func LACM1HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	LACM1HM_func LACM1HM_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D);


	buf MGM_G1(ENABLE_D,D);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACM2HM( Q, QB, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACM2HM_func LACM2HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	LACM2HM_func LACM2HM_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D);


	buf MGM_G1(ENABLE_D,D);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 


   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACM4HM( Q, QB, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACM4HM_func LACM4HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	LACM4HM_func LACM4HM_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D);


	buf MGM_G1(ENABLE_D,D);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQM0HM( Q, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQM0HM_func LACQM0HM_behav_inst(.Q(Q),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	LACQM0HM_func LACQM0HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQM1HM( Q, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQM1HM_func LACQM1HM_behav_inst(.Q(Q),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	LACQM1HM_func LACQM1HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQM2HM( Q, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQM2HM_func LACQM2HM_behav_inst(.Q(Q),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	LACQM2HM_func LACQM2HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQM4HM( Q, D, GB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQM4HM_func LACQM4HM_behav_inst(.Q(Q),.D(D),.GB(GB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	LACQM4HM_func LACQM4HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQRSM0HM( Q, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQRSM0HM_func LACQRSM0HM_behav_inst(.Q(Q),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACQRSM0HM_func LACQRSM0HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQRSM1HM( Q, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQRSM1HM_func LACQRSM1HM_behav_inst(.Q(Q),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACQRSM1HM_func LACQRSM1HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQRSM2HM( Q, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQRSM2HM_func LACQRSM2HM_behav_inst(.Q(Q),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACQRSM2HM_func LACQRSM2HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACQRSM4HM( Q, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACQRSM4HM_func LACQRSM4HM_behav_inst(.Q(Q),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACQRSM4HM_func LACQRSM4HM_inst(.Q(Q),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACRSM0HM( Q, QB, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACRSM0HM_func LACRSM0HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACRSM0HM_func LACRSM0HM_inst(.Q(Q),.QB(QB),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACRSM1HM( Q, QB, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACRSM1HM_func LACRSM1HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACRSM1HM_func LACRSM1HM_inst(.Q(Q),.QB(QB),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACRSM2HM( Q, QB, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACRSM2HM_func LACRSM2HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACRSM2HM_func LACRSM2HM_inst(.Q(Q),.QB(QB),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LACRSM4HM( Q, QB, D, GB, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LACRSM4HM_func LACRSM4HM_behav_inst(.Q(Q),.QB(QB),.D(D),.GB(GB),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire GB$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LACRSM4HM_func LACRSM4HM_inst(.Q(Q),.QB(QB),.D(D$delay),.GB(GB$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	and MGM_G8(MGM_W4,GB$delay,MGM_W3);


	and MGM_G9(ENABLE_NOT_D_AND_GB_AND_SB,SB$delay,MGM_W4);


	and MGM_G10(MGM_W5,GB$delay,D$delay);


	and MGM_G11(ENABLE_D_AND_GB_AND_SB,SB$delay,MGM_W5);


	buf MGM_G12(ENABLE_RB,RB$delay);


	not MGM_G13(MGM_W6,D$delay);


	and MGM_G14(ENABLE_NOT_D_AND_GB,GB$delay,MGM_W6);


	and MGM_G15(ENABLE_D_AND_GB,GB$delay,D$delay);


	not MGM_G16(MGM_W7,D$delay);


	and MGM_G17(MGM_W8,GB$delay,MGM_W7);


	and MGM_G18(ENABLE_NOT_D_AND_GB_AND_RB,RB$delay,MGM_W8);


	and MGM_G19(MGM_W9,GB$delay,D$delay);


	and MGM_G20(ENABLE_D_AND_GB_AND_RB,RB$delay,MGM_W9);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge GB &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_GB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_GB === 1'b1),
		posedge SB &&& (ENABLE_D_AND_GB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_GB_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw GB_hl 
	$width(negedge GB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM12HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM12HM_func LAGCECSM12HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM12HM_func LAGCECSM12HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM16HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM16HM_func LAGCECSM16HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM16HM_func LAGCECSM16HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM20HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM20HM_func LAGCECSM20HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM20HM_func LAGCECSM20HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM2HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM2HM_func LAGCECSM2HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM2HM_func LAGCECSM2HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM3HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM3HM_func LAGCECSM3HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM3HM_func LAGCECSM3HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM4HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM4HM_func LAGCECSM4HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM4HM_func LAGCECSM4HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM6HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM6HM_func LAGCECSM6HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM6HM_func LAGCECSM6HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCECSM8HM( GCK, CKB, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM8HM_func LAGCECSM8HM_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM8HM_func LAGCECSM8HM_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM12HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM12HM_func LAGCEM12HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM12HM_func LAGCEM12HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM16HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM16HM_func LAGCEM16HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM16HM_func LAGCEM16HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM20HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM20HM_func LAGCEM20HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM20HM_func LAGCEM20HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM2HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM2HM_func LAGCEM2HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM2HM_func LAGCEM2HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM3HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM3HM_func LAGCEM3HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM3HM_func LAGCEM3HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM4HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM4HM_func LAGCEM4HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM4HM_func LAGCEM4HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM6HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM6HM_func LAGCEM6HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM6HM_func LAGCEM6HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCEM8HM( GCK, CK, E, VDD, VSS);
inout VDD;
inout VSS;
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM8HM_func LAGCEM8HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM8HM_func LAGCEM8HM_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(ENABLE_NOT_E,E$delay);


	buf MGM_AG1(ENABLE_E,E$delay);


// specify block begins

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM12HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM12HM_func LAGCESM12HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM12HM_func LAGCESM12HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM16HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM16HM_func LAGCESM16HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM16HM_func LAGCESM16HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM20HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM20HM_func LAGCESM20HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM20HM_func LAGCESM20HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM2HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM2HM_func LAGCESM2HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM2HM_func LAGCESM2HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM3HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM3HM_func LAGCESM3HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM3HM_func LAGCESM3HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM4HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM4HM_func LAGCESM4HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM4HM_func LAGCESM4HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM6HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM6HM_func LAGCESM6HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM6HM_func LAGCESM6HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAGCESM8HM( GCK, CK, E, SE, VDD, VSS);
inout VDD;
inout VSS;
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM8HM_func LAGCESM8HM_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM8HM_func LAGCESM8HM_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


	// spec_gates_begin


	not MGM_AG0(MGM_W0,E$delay);


	not MGM_AG1(MGM_W1,SE$delay);


	and MGM_AG2(ENABLE_NOT_E_AND_NOT_SE,MGM_W1,MGM_W0);


	not MGM_AG3(MGM_W2,E$delay);


	and MGM_AG4(ENABLE_NOT_E_AND_SE,SE$delay,MGM_W2);


	not MGM_AG5(MGM_W3,SE$delay);


	and MGM_AG6(ENABLE_E_AND_NOT_SE,MGM_W3,E$delay);


	and MGM_AG7(ENABLE_E_AND_SE,SE$delay,E$delay);


// specify block begins

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_NOT_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK &&& (ENABLE_E_AND_SE === 1'b1)
		,1.0,0,notifier);
	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAM0HM( Q, QB, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAM0HM_func LAM0HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAM0HM_func LAM0HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAM1HM( Q, QB, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAM1HM_func LAM1HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAM1HM_func LAM1HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAM2HM( Q, QB, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAM2HM_func LAM2HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAM2HM_func LAM2HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAM4HM( Q, QB, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAM4HM_func LAM4HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAM4HM_func LAM4HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQM0HM( Q, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQM0HM_func LAQM0HM_behav_inst(.Q(Q),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAQM0HM_func LAQM0HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQM1HM( Q, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQM1HM_func LAQM1HM_behav_inst(.Q(Q),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAQM1HM_func LAQM1HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQM2HM( Q, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQM2HM_func LAQM2HM_behav_inst(.Q(Q),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAQM2HM_func LAQM2HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQM4HM( Q, D, G , VDD, VSS);
inout VDD;
inout VSS;
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQM4HM_func LAQM4HM_behav_inst(.Q(Q),.D(D),.G(G),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	LAQM4HM_func LAQM4HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(ENABLE_NOT_D,D$delay);


	buf MGM_G1(ENABLE_D,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQRSM0HM( Q, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQRSM0HM_func LAQRSM0HM_behav_inst(.Q(Q),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LAQRSM0HM_func LAQRSM0HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQRSM1HM( Q, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQRSM1HM_func LAQRSM1HM_behav_inst(.Q(Q),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LAQRSM1HM_func LAQRSM1HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQRSM2HM( Q, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQRSM2HM_func LAQRSM2HM_behav_inst(.Q(Q),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LAQRSM2HM_func LAQRSM2HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LAQRSM4HM( Q, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LAQRSM4HM_func LAQRSM4HM_behav_inst(.Q(Q),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LAQRSM4HM_func LAQRSM4HM_inst(.Q(Q),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LARSM0HM( Q, QB, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LARSM0HM_func LARSM0HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LARSM0HM_func LARSM0HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LARSM1HM( Q, QB, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LARSM1HM_func LARSM1HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LARSM1HM_func LARSM1HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LARSM2HM( Q, QB, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LARSM2HM_func LARSM2HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LARSM2HM_func LARSM2HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module LARSM4HM( Q, QB, D, G, RB, SB , VDD, VSS);
inout VDD;
inout VSS;
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	LARSM4HM_func LARSM4HM_behav_inst(.Q(Q),.QB(QB),.D(D),.G(G),.RB(RB),.SB(SB),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire D$delay ;

	wire G$delay ;

	wire RB$delay ;

	wire SB$delay ;

	LARSM4HM_func LARSM4HM_inst(.Q(Q),.QB(QB),.D(D$delay),.G(G$delay),.RB(RB$delay),.SB(SB$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	and MGM_G0(ENABLE_RB_AND_SB,SB$delay,RB$delay);


	not MGM_G1(MGM_W0,D$delay);


	and MGM_G2(MGM_W1,RB$delay,MGM_W0);


	and MGM_G3(ENABLE_NOT_D_AND_RB_AND_SB,SB$delay,MGM_W1);


	and MGM_G4(MGM_W2,RB$delay,D$delay);


	and MGM_G5(ENABLE_D_AND_RB_AND_SB,SB$delay,MGM_W2);


	buf MGM_G6(ENABLE_SB,SB$delay);


	not MGM_G7(MGM_W3,D$delay);


	not MGM_G8(MGM_W4,G$delay);


	and MGM_G9(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_G_AND_SB,SB$delay,MGM_W5);


	not MGM_G11(MGM_W6,G$delay);


	and MGM_G12(MGM_W7,MGM_W6,D$delay);


	and MGM_G13(ENABLE_D_AND_NOT_G_AND_SB,SB$delay,MGM_W7);


	buf MGM_G14(ENABLE_RB,RB$delay);


	not MGM_G15(MGM_W8,D$delay);


	not MGM_G16(MGM_W9,G$delay);


	and MGM_G17(ENABLE_NOT_D_AND_NOT_G,MGM_W9,MGM_W8);


	not MGM_G18(MGM_W10,G$delay);


	and MGM_G19(ENABLE_D_AND_NOT_G,MGM_W10,D$delay);


	not MGM_G20(MGM_W11,D$delay);


	not MGM_G21(MGM_W12,G$delay);


	and MGM_G22(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_G_AND_RB,RB$delay,MGM_W13);


	not MGM_G24(MGM_W14,G$delay);


	and MGM_G25(MGM_W15,MGM_W14,D$delay);


	and MGM_G26(ENABLE_D_AND_NOT_G_AND_RB,RB$delay,MGM_W15);


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc D --> Q
	 (D => Q) = (1.0,1.0);

	// seq arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// comb arc D --> QB
	 (D => QB) = (1.0,1.0);

	// seq arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G &&& (ENABLE_NOT_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(posedge G &&& (ENABLE_D_AND_RB_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB &&& (ENABLE_NOT_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_D_AND_NOT_G_AND_SB === 1'b1)
		,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_D_AND_NOT_G === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_D_AND_NOT_G_AND_RB === 1'b1)
		,1.0,0,notifier);

	// mpw G_lh 
	$width(posedge G,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAO222M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAO222M0HM_func MAO222M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAO222M0HM_func MAO222M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAO222M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAO222M1HM_func MAO222M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAO222M1HM_func MAO222M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAO222M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAO222M2HM_func MAO222M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAO222M2HM_func MAO222M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAO222M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAO222M4HM_func MAO222M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAO222M4HM_func MAO222M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI2223M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M0HM_func MAOI2223M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	MAOI2223M0HM_func MAOI2223M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI2223M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M1HM_func MAOI2223M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	MAOI2223M1HM_func MAOI2223M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI2223M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M2HM_func MAOI2223M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	MAOI2223M2HM_func MAOI2223M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI2223M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M4HM_func MAOI2223M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	MAOI2223M4HM_func MAOI2223M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI222M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI222M0HM_func MAOI222M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAOI222M0HM_func MAOI222M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI222M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI222M1HM_func MAOI222M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAOI222M1HM_func MAOI222M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI222M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI222M2HM_func MAOI222M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAOI222M2HM_func MAOI222M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI222M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI222M4HM_func MAOI222M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	MAOI222M4HM_func MAOI222M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI22M0HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI22M0HM_func MAOI22M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MAOI22M0HM_func MAOI22M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI22M1HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI22M1HM_func MAOI22M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MAOI22M1HM_func MAOI22M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI22M2HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI22M2HM_func MAOI22M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MAOI22M2HM_func MAOI22M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MAOI22M4HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MAOI22M4HM_func MAOI22M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MAOI22M4HM_func MAOI22M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MOAI22M0HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MOAI22M0HM_func MOAI22M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MOAI22M0HM_func MOAI22M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MOAI22M1HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MOAI22M1HM_func MOAI22M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MOAI22M1HM_func MOAI22M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MOAI22M2HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MOAI22M2HM_func MOAI22M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MOAI22M2HM_func MOAI22M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MOAI22M4HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MOAI22M4HM_func MOAI22M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	MOAI22M4HM_func MOAI22M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M0HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M0HM_func MUX2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M0HM_func MUX2M0HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M1HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M1HM_func MUX2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M1HM_func MUX2M1HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M2HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M2HM_func MUX2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M2HM_func MUX2M2HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M3HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M3HM_func MUX2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M3HM_func MUX2M3HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M4HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M4HM_func MUX2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M4HM_func MUX2M4HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M6HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M6HM_func MUX2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M6HM_func MUX2M6HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX2M8HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX2M8HM_func MUX2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MUX2M8HM_func MUX2M8HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX3M0HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX3M0HM_func MUX3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX3M0HM_func MUX3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX3M1HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX3M1HM_func MUX3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX3M1HM_func MUX3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX3M2HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX3M2HM_func MUX3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX3M2HM_func MUX3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX3M4HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX3M4HM_func MUX3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX3M4HM_func MUX3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX4M0HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX4M0HM_func MUX4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX4M0HM_func MUX4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX4M1HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX4M1HM_func MUX4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX4M1HM_func MUX4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX4M2HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX4M2HM_func MUX4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX4M2HM_func MUX4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MUX4M4HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MUX4M4HM_func MUX4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MUX4M4HM_func MUX4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M0HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M0HM_func MXB2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M0HM_func MXB2M0HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M1HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M1HM_func MXB2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M1HM_func MXB2M1HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M2HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M2HM_func MXB2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M2HM_func MXB2M2HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M3HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M3HM_func MXB2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M3HM_func MXB2M3HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M4HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M4HM_func MXB2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M4HM_func MXB2M4HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M6HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M6HM_func MXB2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M6HM_func MXB2M6HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB2M8HM( Z, A, B, S , VDD, VSS);
inout VDD;
inout VSS;
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB2M8HM_func MXB2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));

   `else

	MXB2M8HM_func MXB2M8HM_inst(.Z(Z),.A(A),.B(B),.S(S),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	ifnone
	// comb arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB3M0HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB3M0HM_func MXB3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB3M0HM_func MXB3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB3M1HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB3M1HM_func MXB3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB3M1HM_func MXB3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB3M2HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB3M2HM_func MXB3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB3M2HM_func MXB3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB3M4HM( Z, A, B, C, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB3M4HM_func MXB3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB3M4HM_func MXB3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB4M0HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB4M0HM_func MXB4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB4M0HM_func MXB4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB4M1HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB4M1HM_func MXB4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB4M1HM_func MXB4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB4M2HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB4M2HM_func MXB4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB4M2HM_func MXB4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module MXB4M4HM( Z, A, B, C, D, S0, S1 , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	MXB4M4HM_func MXB4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));

   `else

	MXB4M4HM_func MXB4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	ifnone
	// comb arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// comb arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

	ifnone
	// comb arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// comb arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2B1M0HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2B1M0HM_func ND2B1M0HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND2B1M0HM_func ND2B1M0HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2B1M12HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2B1M12HM_func ND2B1M12HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND2B1M12HM_func ND2B1M12HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2B1M1HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2B1M1HM_func ND2B1M1HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND2B1M1HM_func ND2B1M1HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2B1M2HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2B1M2HM_func ND2B1M2HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND2B1M2HM_func ND2B1M2HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2B1M4HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2B1M4HM_func ND2B1M4HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND2B1M4HM_func ND2B1M4HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2B1M8HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2B1M8HM_func ND2B1M8HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND2B1M8HM_func ND2B1M8HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M0HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M0HM_func ND2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M0HM_func ND2M0HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M12HM_func ND2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M12HM_func ND2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M16HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M16HM_func ND2M16HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M16HM_func ND2M16HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M1HM_func ND2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M1HM_func ND2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M2HM_func ND2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M2HM_func ND2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M3HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M3HM_func ND2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M3HM_func ND2M3HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M4HM_func ND2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M4HM_func ND2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M5HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M5HM_func ND2M5HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M5HM_func ND2M5HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M6HM_func ND2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M6HM_func ND2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND2M8HM_func ND2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	ND2M8HM_func ND2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3B1M0HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3B1M0HM_func ND3B1M0HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND3B1M0HM_func ND3B1M0HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3B1M1HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3B1M1HM_func ND3B1M1HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND3B1M1HM_func ND3B1M1HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3B1M2HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3B1M2HM_func ND3B1M2HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND3B1M2HM_func ND3B1M2HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3B1M4HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3B1M4HM_func ND3B1M4HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND3B1M4HM_func ND3B1M4HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3B1M8HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3B1M8HM_func ND3B1M8HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND3B1M8HM_func ND3B1M8HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M0HM_func ND3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M0HM_func ND3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M12HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M12HM_func ND3M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M12HM_func ND3M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M16HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M16HM_func ND3M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M16HM_func ND3M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M1HM_func ND3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M1HM_func ND3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M2HM_func ND3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M2HM_func ND3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M3HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M3HM_func ND3M3HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M3HM_func ND3M3HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M4HM_func ND3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M4HM_func ND3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M6HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M6HM_func ND3M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M6HM_func ND3M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND3M8HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND3M8HM_func ND3M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	ND3M8HM_func ND3M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B1M0HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B1M0HM_func ND4B1M0HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND4B1M0HM_func ND4B1M0HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B1M1HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B1M1HM_func ND4B1M1HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND4B1M1HM_func ND4B1M1HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B1M2HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B1M2HM_func ND4B1M2HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND4B1M2HM_func ND4B1M2HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B1M4HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B1M4HM_func ND4B1M4HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND4B1M4HM_func ND4B1M4HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B1M8HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B1M8HM_func ND4B1M8HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	ND4B1M8HM_func ND4B1M8HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B2M0HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B2M0HM_func ND4B2M0HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	ND4B2M0HM_func ND4B2M0HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B2M1HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B2M1HM_func ND4B2M1HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	ND4B2M1HM_func ND4B2M1HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B2M2HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B2M2HM_func ND4B2M2HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	ND4B2M2HM_func ND4B2M2HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B2M4HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B2M4HM_func ND4B2M4HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	ND4B2M4HM_func ND4B2M4HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4B2M8HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4B2M8HM_func ND4B2M8HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	ND4B2M8HM_func ND4B2M8HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M0HM_func ND4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M0HM_func ND4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M12HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M12HM_func ND4M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M12HM_func ND4M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M16HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M16HM_func ND4M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M16HM_func ND4M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M1HM_func ND4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M1HM_func ND4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M2HM_func ND4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M2HM_func ND4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M4HM_func ND4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M4HM_func ND4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M6HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M6HM_func ND4M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M6HM_func ND4M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ND4M8HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	ND4M8HM_func ND4M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	ND4M8HM_func ND4M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2B1M0HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2B1M0HM_func NR2B1M0HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR2B1M0HM_func NR2B1M0HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2B1M12HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2B1M12HM_func NR2B1M12HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR2B1M12HM_func NR2B1M12HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2B1M1HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2B1M1HM_func NR2B1M1HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR2B1M1HM_func NR2B1M1HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2B1M2HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2B1M2HM_func NR2B1M2HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR2B1M2HM_func NR2B1M2HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2B1M4HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2B1M4HM_func NR2B1M4HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR2B1M4HM_func NR2B1M4HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2B1M8HM( Z, B, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2B1M8HM_func NR2B1M8HM_behav_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR2B1M8HM_func NR2B1M8HM_inst(.Z(Z),.B(B),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M0HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M0HM_func NR2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M0HM_func NR2M0HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M12HM_func NR2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M12HM_func NR2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M16HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M16HM_func NR2M16HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M16HM_func NR2M16HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M1HM_func NR2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M1HM_func NR2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M2HM_func NR2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M2HM_func NR2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M3HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M3HM_func NR2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M3HM_func NR2M3HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M4HM_func NR2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M4HM_func NR2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M5HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M5HM_func NR2M5HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M5HM_func NR2M5HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M6HM_func NR2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M6HM_func NR2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR2M8HM_func NR2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	NR2M8HM_func NR2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3B1M0HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3B1M0HM_func NR3B1M0HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR3B1M0HM_func NR3B1M0HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3B1M1HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3B1M1HM_func NR3B1M1HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR3B1M1HM_func NR3B1M1HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3B1M2HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3B1M2HM_func NR3B1M2HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR3B1M2HM_func NR3B1M2HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3B1M4HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3B1M4HM_func NR3B1M4HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR3B1M4HM_func NR3B1M4HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3B1M8HM( Z, B, C, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3B1M8HM_func NR3B1M8HM_behav_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR3B1M8HM_func NR3B1M8HM_inst(.Z(Z),.B(B),.C(C),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M0HM_func NR3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M0HM_func NR3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M12HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M12HM_func NR3M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M12HM_func NR3M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M16HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M16HM_func NR3M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M16HM_func NR3M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M1HM_func NR3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M1HM_func NR3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M2HM_func NR3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M2HM_func NR3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M4HM_func NR3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M4HM_func NR3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M6HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M6HM_func NR3M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M6HM_func NR3M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR3M8HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR3M8HM_func NR3M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	NR3M8HM_func NR3M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B1M0HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B1M0HM_func NR4B1M0HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR4B1M0HM_func NR4B1M0HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B1M1HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B1M1HM_func NR4B1M1HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR4B1M1HM_func NR4B1M1HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B1M2HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B1M2HM_func NR4B1M2HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR4B1M2HM_func NR4B1M2HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B1M4HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B1M4HM_func NR4B1M4HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR4B1M4HM_func NR4B1M4HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B1M8HM( Z, B, C, D, NA , VDD, VSS);
inout VDD;
inout VSS;
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B1M8HM_func NR4B1M8HM_behav_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));

   `else

	NR4B1M8HM_func NR4B1M8HM_inst(.Z(Z),.B(B),.C(C),.D(D),.NA(NA),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B2M0HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B2M0HM_func NR4B2M0HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	NR4B2M0HM_func NR4B2M0HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B2M1HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B2M1HM_func NR4B2M1HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	NR4B2M1HM_func NR4B2M1HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B2M2HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B2M2HM_func NR4B2M2HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	NR4B2M2HM_func NR4B2M2HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B2M4HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B2M4HM_func NR4B2M4HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	NR4B2M4HM_func NR4B2M4HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4B2M8HM( Z, C, D, NA, NB , VDD, VSS);
inout VDD;
inout VSS;
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4B2M8HM_func NR4B2M8HM_behav_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	NR4B2M8HM_func NR4B2M8HM_inst(.Z(Z),.C(C),.D(D),.NA(NA),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M0HM_func NR4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M0HM_func NR4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M12HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M12HM_func NR4M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M12HM_func NR4M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M16HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M16HM_func NR4M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M16HM_func NR4M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M1HM_func NR4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M1HM_func NR4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M2HM_func NR4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M2HM_func NR4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M4HM_func NR4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M4HM_func NR4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M6HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M6HM_func NR4M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M6HM_func NR4M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module NR4M8HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	NR4M8HM_func NR4M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	NR4M8HM_func NR4M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA211M0HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA211M0HM_func OA211M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA211M0HM_func OA211M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA211M1HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA211M1HM_func OA211M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA211M1HM_func OA211M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA211M2HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA211M2HM_func OA211M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA211M2HM_func OA211M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA211M4HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA211M4HM_func OA211M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA211M4HM_func OA211M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA211M8HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA211M8HM_func OA211M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA211M8HM_func OA211M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA21M0HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA21M0HM_func OA21M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA21M0HM_func OA21M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA21M1HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA21M1HM_func OA21M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA21M1HM_func OA21M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA21M2HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA21M2HM_func OA21M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA21M2HM_func OA21M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA21M4HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA21M4HM_func OA21M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA21M4HM_func OA21M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA21M8HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA21M8HM_func OA21M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA21M8HM_func OA21M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA221M0HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA221M0HM_func OA221M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA221M0HM_func OA221M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA221M1HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA221M1HM_func OA221M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA221M1HM_func OA221M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA221M2HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA221M2HM_func OA221M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA221M2HM_func OA221M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA221M4HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA221M4HM_func OA221M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA221M4HM_func OA221M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA221M8HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA221M8HM_func OA221M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OA221M8HM_func OA221M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA222M0HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA222M0HM_func OA222M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OA222M0HM_func OA222M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA222M1HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA222M1HM_func OA222M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OA222M1HM_func OA222M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA222M2HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA222M2HM_func OA222M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OA222M2HM_func OA222M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA222M4HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA222M4HM_func OA222M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OA222M4HM_func OA222M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA222M8HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA222M8HM_func OA222M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OA222M8HM_func OA222M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA22M0HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA22M0HM_func OA22M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA22M0HM_func OA22M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA22M1HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA22M1HM_func OA22M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA22M1HM_func OA22M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA22M2HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA22M2HM_func OA22M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA22M2HM_func OA22M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA22M4HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA22M4HM_func OA22M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA22M4HM_func OA22M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA22M8HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA22M8HM_func OA22M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA22M8HM_func OA22M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA31M0HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA31M0HM_func OA31M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA31M0HM_func OA31M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA31M1HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA31M1HM_func OA31M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA31M1HM_func OA31M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA31M2HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA31M2HM_func OA31M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA31M2HM_func OA31M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA31M4HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA31M4HM_func OA31M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA31M4HM_func OA31M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA31M8HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA31M8HM_func OA31M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OA31M8HM_func OA31M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA32M0HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA32M0HM_func OA32M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA32M0HM_func OA32M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA32M1HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA32M1HM_func OA32M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA32M1HM_func OA32M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA32M2HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA32M2HM_func OA32M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA32M2HM_func OA32M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA32M4HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA32M4HM_func OA32M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA32M4HM_func OA32M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA32M8HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA32M8HM_func OA32M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OA32M8HM_func OA32M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA33M0HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA33M0HM_func OA33M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OA33M0HM_func OA33M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA33M1HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA33M1HM_func OA33M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OA33M1HM_func OA33M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA33M2HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA33M2HM_func OA33M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OA33M2HM_func OA33M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA33M4HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA33M4HM_func OA33M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OA33M4HM_func OA33M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OA33M8HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OA33M8HM_func OA33M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OA33M8HM_func OA33M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211B100M0HM( Z, A1, B, C, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M0HM_func OAI211B100M0HM_behav_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI211B100M0HM_func OAI211B100M0HM_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211B100M1HM( Z, A1, B, C, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M1HM_func OAI211B100M1HM_behav_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI211B100M1HM_func OAI211B100M1HM_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211B100M2HM( Z, A1, B, C, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M2HM_func OAI211B100M2HM_behav_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI211B100M2HM_func OAI211B100M2HM_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211B100M4HM( Z, A1, B, C, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M4HM_func OAI211B100M4HM_behav_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI211B100M4HM_func OAI211B100M4HM_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211B100M8HM( Z, A1, B, C, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M8HM_func OAI211B100M8HM_behav_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI211B100M8HM_func OAI211B100M8HM_inst(.Z(Z),.A1(A1),.B(B),.C(C),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211M0HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211M0HM_func OAI211M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI211M0HM_func OAI211M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211M1HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211M1HM_func OAI211M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI211M1HM_func OAI211M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211M2HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211M2HM_func OAI211M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI211M2HM_func OAI211M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211M4HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211M4HM_func OAI211M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI211M4HM_func OAI211M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI211M8HM( Z, A1, A2, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI211M8HM_func OAI211M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI211M8HM_func OAI211M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B01M0HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M0HM_func OAI21B01M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B01M0HM_func OAI21B01M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B01M1HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M1HM_func OAI21B01M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B01M1HM_func OAI21B01M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B01M2HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M2HM_func OAI21B01M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B01M2HM_func OAI21B01M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B01M4HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M4HM_func OAI21B01M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B01M4HM_func OAI21B01M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B01M8HM( Z, A1, A2, NB , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M8HM_func OAI21B01M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B01M8HM_func OAI21B01M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.NB(NB),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// comb arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B10M0HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M0HM_func OAI21B10M0HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B10M0HM_func OAI21B10M0HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B10M1HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M1HM_func OAI21B10M1HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B10M1HM_func OAI21B10M1HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B10M2HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M2HM_func OAI21B10M2HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B10M2HM_func OAI21B10M2HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B10M4HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M4HM_func OAI21B10M4HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B10M4HM_func OAI21B10M4HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B10M8HM( Z, A1, B, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M8HM_func OAI21B10M8HM_behav_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B10M8HM_func OAI21B10M8HM_inst(.Z(Z),.A1(A1),.B(B),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B20M0HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M0HM_func OAI21B20M0HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B20M0HM_func OAI21B20M0HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B20M1HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M1HM_func OAI21B20M1HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B20M1HM_func OAI21B20M1HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B20M2HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M2HM_func OAI21B20M2HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B20M2HM_func OAI21B20M2HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B20M4HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M4HM_func OAI21B20M4HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B20M4HM_func OAI21B20M4HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21B20M8HM( Z, B, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M8HM_func OAI21B20M8HM_behav_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI21B20M8HM_func OAI21B20M8HM_inst(.Z(Z),.B(B),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M0HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M0HM_func OAI21M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M0HM_func OAI21M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M1HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M1HM_func OAI21M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M1HM_func OAI21M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M2HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M2HM_func OAI21M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M2HM_func OAI21M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M3HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M3HM_func OAI21M3HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M3HM_func OAI21M3HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M4HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M4HM_func OAI21M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M4HM_func OAI21M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M6HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M6HM_func OAI21M6HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M6HM_func OAI21M6HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI21M8HM( Z, A1, A2, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI21M8HM_func OAI21M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI21M8HM_func OAI21M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI221M0HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI221M0HM_func OAI221M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI221M0HM_func OAI221M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI221M1HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI221M1HM_func OAI221M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI221M1HM_func OAI221M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI221M2HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI221M2HM_func OAI221M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI221M2HM_func OAI221M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI221M4HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI221M4HM_func OAI221M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI221M4HM_func OAI221M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI221M8HM( Z, A1, A2, B1, B2, C , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI221M8HM_func OAI221M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OAI221M8HM_func OAI221M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI222M0HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI222M0HM_func OAI222M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OAI222M0HM_func OAI222M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI222M1HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI222M1HM_func OAI222M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OAI222M1HM_func OAI222M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI222M2HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI222M2HM_func OAI222M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OAI222M2HM_func OAI222M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI222M4HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI222M4HM_func OAI222M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OAI222M4HM_func OAI222M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI222M8HM( Z, A1, A2, B1, B2, C1, C2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI222M8HM_func OAI222M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));

   `else

	OAI222M8HM_func OAI222M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// comb arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// comb arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B10M0HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M0HM_func OAI22B10M0HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B10M0HM_func OAI22B10M0HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B10M1HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M1HM_func OAI22B10M1HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B10M1HM_func OAI22B10M1HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B10M2HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M2HM_func OAI22B10M2HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B10M2HM_func OAI22B10M2HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B10M4HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M4HM_func OAI22B10M4HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B10M4HM_func OAI22B10M4HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B10M8HM( Z, A1, B1, B2, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M8HM_func OAI22B10M8HM_behav_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B10M8HM_func OAI22B10M8HM_inst(.Z(Z),.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B20M0HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M0HM_func OAI22B20M0HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B20M0HM_func OAI22B20M0HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B20M1HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M1HM_func OAI22B20M1HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B20M1HM_func OAI22B20M1HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B20M2HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M2HM_func OAI22B20M2HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B20M2HM_func OAI22B20M2HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B20M4HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M4HM_func OAI22B20M4HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B20M4HM_func OAI22B20M4HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22B20M8HM( Z, B1, B2, NA1, NA2 , VDD, VSS);
inout VDD;
inout VSS;
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M8HM_func OAI22B20M8HM_behav_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22B20M8HM_func OAI22B20M8HM_inst(.Z(Z),.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// comb arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22M0HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22M0HM_func OAI22M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22M0HM_func OAI22M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22M1HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22M1HM_func OAI22M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22M1HM_func OAI22M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22M2HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22M2HM_func OAI22M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22M2HM_func OAI22M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22M4HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22M4HM_func OAI22M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22M4HM_func OAI22M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI22M8HM( Z, A1, A2, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI22M8HM_func OAI22M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI22M8HM_func OAI22M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI31M0HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI31M0HM_func OAI31M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI31M0HM_func OAI31M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI31M1HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI31M1HM_func OAI31M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI31M1HM_func OAI31M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI31M2HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI31M2HM_func OAI31M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI31M2HM_func OAI31M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI31M4HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI31M4HM_func OAI31M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI31M4HM_func OAI31M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI31M8HM( Z, A1, A2, A3, B , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI31M8HM_func OAI31M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OAI31M8HM_func OAI31M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI32M0HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI32M0HM_func OAI32M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI32M0HM_func OAI32M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI32M1HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI32M1HM_func OAI32M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI32M1HM_func OAI32M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI32M2HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI32M2HM_func OAI32M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI32M2HM_func OAI32M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI32M4HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI32M4HM_func OAI32M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI32M4HM_func OAI32M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI32M8HM( Z, A1, A2, A3, B1, B2 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI32M8HM_func OAI32M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));

   `else

	OAI32M8HM_func OAI32M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI33M0HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI33M0HM_func OAI33M0HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OAI33M0HM_func OAI33M0HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI33M1HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI33M1HM_func OAI33M1HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OAI33M1HM_func OAI33M1HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI33M2HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI33M2HM_func OAI33M2HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OAI33M2HM_func OAI33M2HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI33M4HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI33M4HM_func OAI33M4HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OAI33M4HM_func OAI33M4HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OAI33M8HM( Z, A1, A2, A3, B1, B2, B3 , VDD, VSS);
inout VDD;
inout VSS;
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OAI33M8HM_func OAI33M8HM_behav_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));

   `else

	OAI33M8HM_func OAI33M8HM_inst(.Z(Z),.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// comb arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// comb arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// comb arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// comb arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// comb arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// comb arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M0HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M0HM_func OR2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M0HM_func OR2M0HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M12HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M12HM_func OR2M12HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M12HM_func OR2M12HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M16HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M16HM_func OR2M16HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M16HM_func OR2M16HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M1HM_func OR2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M1HM_func OR2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M2HM_func OR2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M2HM_func OR2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M4HM_func OR2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M4HM_func OR2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M6HM_func OR2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M6HM_func OR2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR2M8HM_func OR2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	OR2M8HM_func OR2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M0HM_func OR3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M0HM_func OR3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M12HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M12HM_func OR3M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M12HM_func OR3M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M16HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M16HM_func OR3M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M16HM_func OR3M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M1HM_func OR3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M1HM_func OR3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M2HM_func OR3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M2HM_func OR3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M4HM_func OR3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M4HM_func OR3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M6HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M6HM_func OR3M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M6HM_func OR3M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR3M8HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR3M8HM_func OR3M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	OR3M8HM_func OR3M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M0HM_func OR4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M0HM_func OR4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M12HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M12HM_func OR4M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M12HM_func OR4M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M16HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M16HM_func OR4M16HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M16HM_func OR4M16HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M1HM_func OR4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M1HM_func OR4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M2HM_func OR4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M2HM_func OR4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M4HM_func OR4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M4HM_func OR4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M6HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M6HM_func OR4M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M6HM_func OR4M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR4M8HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR4M8HM_func OR4M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	OR4M8HM_func OR4M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M0HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M0HM_func OR6M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M0HM_func OR6M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M12HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M12HM_func OR6M12HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M12HM_func OR6M12HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M1HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M1HM_func OR6M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M1HM_func OR6M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M2HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M2HM_func OR6M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M2HM_func OR6M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M4HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M4HM_func OR6M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M4HM_func OR6M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M6HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M6HM_func OR6M6HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M6HM_func OR6M6HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module OR6M8HM( Z, A, B, C, D, E, F , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	OR6M8HM_func OR6M8HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));

   `else

	OR6M8HM_func OR6M8HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// comb arc E --> Z
	 (E => Z) = (1.0,1.0);

	// comb arc F --> Z
	 (F => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCM1HM( Q, QB, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCM1HM_func SDFCM1HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCM1HM_func SDFCM1HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCM2HM( Q, QB, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCM2HM_func SDFCM2HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCM2HM_func SDFCM2HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCM4HM( Q, QB, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCM4HM_func SDFCM4HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCM4HM_func SDFCM4HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCM8HM( Q, QB, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCM8HM_func SDFCM8HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCM8HM_func SDFCM8HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQM1HM( Q, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQM1HM_func SDFCQM1HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQM1HM_func SDFCQM1HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQM2HM( Q, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQM2HM_func SDFCQM2HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQM2HM_func SDFCQM2HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQM4HM( Q, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQM4HM_func SDFCQM4HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQM4HM_func SDFCQM4HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQM8HM( Q, CKB, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQM8HM_func SDFCQM8HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQM8HM_func SDFCQM8HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQRSM1HM( Q, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM1HM_func SDFCQRSM1HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQRSM1HM_func SDFCQRSM1HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQRSM2HM( Q, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM2HM_func SDFCQRSM2HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQRSM2HM_func SDFCQRSM2HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQRSM4HM( Q, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM4HM_func SDFCQRSM4HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQRSM4HM_func SDFCQRSM4HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCQRSM8HM( Q, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM8HM_func SDFCQRSM8HM_behav_inst(.Q(Q),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCQRSM8HM_func SDFCQRSM8HM_inst(.Q(Q),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCRSM1HM( Q, QB, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM1HM_func SDFCRSM1HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCRSM1HM_func SDFCRSM1HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCRSM2HM( Q, QB, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM2HM_func SDFCRSM2HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCRSM2HM_func SDFCRSM2HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCRSM4HM( Q, QB, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM4HM_func SDFCRSM4HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCRSM4HM_func SDFCRSM4HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFCRSM8HM( Q, QB, CKB, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM8HM_func SDFCRSM8HM_behav_inst(.Q(Q),.QB(QB),.CKB(CKB),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CKB$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFCRSM8HM_func SDFCRSM8HM_inst(.Q(Q),.QB(QB),.CKB(CKB$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CKB$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CKB$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CKB$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CKB$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CKB$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CKB$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CKB$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CKB$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CKB$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CKB$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CKB$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CKB$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CKB$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CKB$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CKB$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CKB$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CKB$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CKB$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CKB$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CKB$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CKB$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CKB$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CKB$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CKB$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CKB$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CKB$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CKB$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CKB$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CKB$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CKB$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CKB$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CKB$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CKB_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CKB$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CKB$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CKB$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CKB$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CKB$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CKB$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CKB$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CKB$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CKB$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CKB$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CKB$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CKB$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CKB$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CKB$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CKB$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CKB$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CKB_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		negedge CKB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CKB_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CKB_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// mpw CKB_lh 
	$width(posedge CKB,1.0,0,notifier);

	// mpw CKB_hl 
	$width(negedge CKB,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEM1HM( Q, QB, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEM1HM_func SDFEM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEM1HM_func SDFEM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEM2HM( Q, QB, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEM2HM_func SDFEM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEM2HM_func SDFEM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEM4HM( Q, QB, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEM4HM_func SDFEM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEM4HM_func SDFEM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEM8HM( Q, QB, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEM8HM_func SDFEM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEM8HM_func SDFEM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQM1HM( Q, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQM1HM_func SDFEQM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQM1HM_func SDFEQM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQM2HM( Q, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQM2HM_func SDFEQM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQM2HM_func SDFEQM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQM4HM( Q, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQM4HM_func SDFEQM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQM4HM_func SDFEQM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQM8HM( Q, CK, D, E, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQM8HM_func SDFEQM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQM8HM_func SDFEQM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	and MGM_G5(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W4);


	not MGM_G6(MGM_W5,D$delay);


	not MGM_G7(MGM_W6,E$delay);


	and MGM_G8(MGM_W7,MGM_W6,MGM_W5);


	and MGM_G9(MGM_W8,SD$delay,MGM_W7);


	and MGM_G10(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,E$delay,MGM_W9);


	not MGM_G13(MGM_W11,SD$delay);


	and MGM_G14(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G15(MGM_W13,SE$delay);


	and MGM_G16(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W13,MGM_W12);


	not MGM_G17(MGM_W14,D$delay);


	and MGM_G18(MGM_W15,E$delay,MGM_W14);


	not MGM_G19(MGM_W16,SD$delay);


	and MGM_G20(MGM_W17,MGM_W16,MGM_W15);


	and MGM_G21(ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W17);


	not MGM_G22(MGM_W18,D$delay);


	and MGM_G23(MGM_W19,E$delay,MGM_W18);


	and MGM_G24(MGM_W20,SD$delay,MGM_W19);


	not MGM_G25(MGM_W21,SE$delay);


	and MGM_G26(ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G27(MGM_W22,D$delay);


	and MGM_G28(MGM_W23,E$delay,MGM_W22);


	and MGM_G29(MGM_W24,SD$delay,MGM_W23);


	and MGM_G30(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W24);


	not MGM_G31(MGM_W25,E$delay);


	and MGM_G32(MGM_W26,MGM_W25,D$delay);


	not MGM_G33(MGM_W27,SD$delay);


	and MGM_G34(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G35(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G36(MGM_W29,E$delay);


	and MGM_G37(MGM_W30,MGM_W29,D$delay);


	and MGM_G38(MGM_W31,SD$delay,MGM_W30);


	and MGM_G39(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W31);


	and MGM_G40(MGM_W32,E$delay,D$delay);


	not MGM_G41(MGM_W33,SD$delay);


	and MGM_G42(MGM_W34,MGM_W33,MGM_W32);


	not MGM_G43(MGM_W35,SE$delay);


	and MGM_G44(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W35,MGM_W34);


	and MGM_G45(MGM_W36,E$delay,D$delay);


	not MGM_G46(MGM_W37,SD$delay);


	and MGM_G47(MGM_W38,MGM_W37,MGM_W36);


	and MGM_G48(ENABLE_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W38);


	and MGM_G49(MGM_W39,E$delay,D$delay);


	and MGM_G50(MGM_W40,SD$delay,MGM_W39);


	not MGM_G51(MGM_W41,SE$delay);


	and MGM_G52(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W41,MGM_W40);


	and MGM_G53(MGM_W42,E$delay,D$delay);


	and MGM_G54(MGM_W43,SD$delay,MGM_W42);


	and MGM_G55(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W43);


	not MGM_G56(MGM_W44,SD$delay);


	and MGM_G57(MGM_W45,MGM_W44,E$delay);


	not MGM_G58(MGM_W46,SE$delay);


	and MGM_G59(ENABLE_E_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	and MGM_G60(MGM_W47,SD$delay,E$delay);


	not MGM_G61(MGM_W48,SE$delay);


	and MGM_G62(ENABLE_E_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G63(MGM_W49,D$delay);


	not MGM_G64(MGM_W50,SD$delay);


	and MGM_G65(MGM_W51,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W52,SE$delay);


	and MGM_G67(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	not MGM_G68(MGM_W53,D$delay);


	and MGM_G69(MGM_W54,SD$delay,MGM_W53);


	not MGM_G70(MGM_W55,SE$delay);


	and MGM_G71(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	not MGM_G72(MGM_W56,SD$delay);


	and MGM_G73(MGM_W57,MGM_W56,D$delay);


	not MGM_G74(MGM_W58,SE$delay);


	and MGM_G75(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	and MGM_G76(MGM_W59,SD$delay,D$delay);


	not MGM_G77(MGM_W60,SE$delay);


	and MGM_G78(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G79(MGM_W61,D$delay);


	not MGM_G80(MGM_W62,E$delay);


	and MGM_G81(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G82(ENABLE_NOT_D_AND_NOT_E_AND_SE,SE$delay,MGM_W63);


	not MGM_G83(MGM_W64,D$delay);


	and MGM_G84(MGM_W65,E$delay,MGM_W64);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_SE,SE$delay,MGM_W65);


	not MGM_G86(MGM_W66,E$delay);


	and MGM_G87(MGM_W67,MGM_W66,D$delay);


	and MGM_G88(ENABLE_D_AND_NOT_E_AND_SE,SE$delay,MGM_W67);


	and MGM_G89(MGM_W68,E$delay,D$delay);


	and MGM_G90(ENABLE_D_AND_E_AND_SE,SE$delay,MGM_W68);


	not MGM_G91(MGM_W69,D$delay);


	not MGM_G92(MGM_W70,E$delay);


	and MGM_G93(MGM_W71,MGM_W70,MGM_W69);


	not MGM_G94(MGM_W72,SD$delay);


	and MGM_G95(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD,MGM_W72,MGM_W71);


	not MGM_G96(MGM_W73,D$delay);


	not MGM_G97(MGM_W74,E$delay);


	and MGM_G98(MGM_W75,MGM_W74,MGM_W73);


	and MGM_G99(ENABLE_NOT_D_AND_NOT_E_AND_SD,SD$delay,MGM_W75);


	not MGM_G100(MGM_W76,D$delay);


	and MGM_G101(MGM_W77,E$delay,MGM_W76);


	and MGM_G102(ENABLE_NOT_D_AND_E_AND_SD,SD$delay,MGM_W77);


	not MGM_G103(MGM_W78,E$delay);


	and MGM_G104(MGM_W79,MGM_W78,D$delay);


	not MGM_G105(MGM_W80,SD$delay);


	and MGM_G106(ENABLE_D_AND_NOT_E_AND_NOT_SD,MGM_W80,MGM_W79);


	not MGM_G107(MGM_W81,E$delay);


	and MGM_G108(MGM_W82,MGM_W81,D$delay);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD,SD$delay,MGM_W82);


	and MGM_G110(MGM_W83,E$delay,D$delay);


	not MGM_G111(MGM_W84,SD$delay);


	and MGM_G112(ENABLE_D_AND_E_AND_NOT_SD,MGM_W84,MGM_W83);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQRM1HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM1HM_func SDFEQRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQRM1HM_func SDFEQRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQRM2HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM2HM_func SDFEQRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQRM2HM_func SDFEQRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQRM4HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM4HM_func SDFEQRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQRM4HM_func SDFEQRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQRM8HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM8HM_func SDFEQRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQRM8HM_func SDFEQRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQZRM1HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM1HM_func SDFEQZRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQZRM1HM_func SDFEQZRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQZRM2HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM2HM_func SDFEQZRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQZRM2HM_func SDFEQZRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQZRM4HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM4HM_func SDFEQZRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQZRM4HM_func SDFEQZRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEQZRM8HM( Q, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM8HM_func SDFEQZRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEQZRM8HM_func SDFEQZRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFERM1HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFERM1HM_func SDFERM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFERM1HM_func SDFERM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFERM2HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFERM2HM_func SDFERM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFERM2HM_func SDFERM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFERM4HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFERM4HM_func SDFERM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFERM4HM_func SDFERM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFERM8HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFERM8HM_func SDFERM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFERM8HM_func SDFERM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	and MGM_G3(MGM_W3,RB$delay,MGM_W2);


	not MGM_G4(MGM_W4,SD$delay);


	and MGM_G5(MGM_W5,MGM_W4,MGM_W3);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W5);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,E$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(MGM_W9,RB$delay,MGM_W8);


	and MGM_G11(MGM_W10,SD$delay,MGM_W9);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,E$delay,MGM_W11);


	and MGM_G15(MGM_W13,RB$delay,MGM_W12);


	not MGM_G16(MGM_W14,SD$delay);


	and MGM_G17(MGM_W15,MGM_W14,MGM_W13);


	not MGM_G18(MGM_W16,SE$delay);


	and MGM_G19(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W17,D$delay);


	and MGM_G21(MGM_W18,E$delay,MGM_W17);


	and MGM_G22(MGM_W19,RB$delay,MGM_W18);


	not MGM_G23(MGM_W20,SD$delay);


	and MGM_G24(MGM_W21,MGM_W20,MGM_W19);


	and MGM_G25(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W21);


	not MGM_G26(MGM_W22,D$delay);


	and MGM_G27(MGM_W23,E$delay,MGM_W22);


	and MGM_G28(MGM_W24,RB$delay,MGM_W23);


	and MGM_G29(MGM_W25,SD$delay,MGM_W24);


	not MGM_G30(MGM_W26,SE$delay);


	and MGM_G31(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W26,MGM_W25);


	not MGM_G32(MGM_W27,D$delay);


	and MGM_G33(MGM_W28,E$delay,MGM_W27);


	and MGM_G34(MGM_W29,RB$delay,MGM_W28);


	and MGM_G35(MGM_W30,SD$delay,MGM_W29);


	and MGM_G36(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W30);


	not MGM_G37(MGM_W31,E$delay);


	and MGM_G38(MGM_W32,MGM_W31,D$delay);


	and MGM_G39(MGM_W33,RB$delay,MGM_W32);


	not MGM_G40(MGM_W34,SD$delay);


	and MGM_G41(MGM_W35,MGM_W34,MGM_W33);


	and MGM_G42(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G43(MGM_W36,E$delay);


	and MGM_G44(MGM_W37,MGM_W36,D$delay);


	and MGM_G45(MGM_W38,RB$delay,MGM_W37);


	and MGM_G46(MGM_W39,SD$delay,MGM_W38);


	and MGM_G47(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W39);


	and MGM_G48(MGM_W40,E$delay,D$delay);


	and MGM_G49(MGM_W41,RB$delay,MGM_W40);


	not MGM_G50(MGM_W42,SD$delay);


	and MGM_G51(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G52(MGM_W44,SE$delay);


	and MGM_G53(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W44,MGM_W43);


	and MGM_G54(MGM_W45,E$delay,D$delay);


	and MGM_G55(MGM_W46,RB$delay,MGM_W45);


	not MGM_G56(MGM_W47,SD$delay);


	and MGM_G57(MGM_W48,MGM_W47,MGM_W46);


	and MGM_G58(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W48);


	and MGM_G59(MGM_W49,E$delay,D$delay);


	and MGM_G60(MGM_W50,RB$delay,MGM_W49);


	and MGM_G61(MGM_W51,SD$delay,MGM_W50);


	not MGM_G62(MGM_W52,SE$delay);


	and MGM_G63(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G64(MGM_W53,E$delay,D$delay);


	and MGM_G65(MGM_W54,RB$delay,MGM_W53);


	and MGM_G66(MGM_W55,SD$delay,MGM_W54);


	and MGM_G67(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W55);


	and MGM_G68(MGM_W56,RB$delay,E$delay);


	not MGM_G69(MGM_W57,SD$delay);


	and MGM_G70(MGM_W58,MGM_W57,MGM_W56);


	not MGM_G71(MGM_W59,SE$delay);


	and MGM_G72(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W59,MGM_W58);


	and MGM_G73(MGM_W60,RB$delay,E$delay);


	and MGM_G74(MGM_W61,SD$delay,MGM_W60);


	not MGM_G75(MGM_W62,SE$delay);


	and MGM_G76(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W62,MGM_W61);


	not MGM_G77(MGM_W63,D$delay);


	and MGM_G78(MGM_W64,RB$delay,MGM_W63);


	not MGM_G79(MGM_W65,SD$delay);


	and MGM_G80(MGM_W66,MGM_W65,MGM_W64);


	not MGM_G81(MGM_W67,SE$delay);


	and MGM_G82(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W67,MGM_W66);


	not MGM_G83(MGM_W68,D$delay);


	and MGM_G84(MGM_W69,RB$delay,MGM_W68);


	and MGM_G85(MGM_W70,SD$delay,MGM_W69);


	not MGM_G86(MGM_W71,SE$delay);


	and MGM_G87(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G88(MGM_W72,RB$delay,D$delay);


	not MGM_G89(MGM_W73,SD$delay);


	and MGM_G90(MGM_W74,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W75,SE$delay);


	and MGM_G92(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W75,MGM_W74);


	and MGM_G93(MGM_W76,RB$delay,D$delay);


	and MGM_G94(MGM_W77,SD$delay,MGM_W76);


	not MGM_G95(MGM_W78,SE$delay);


	and MGM_G96(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G97(MGM_W79,D$delay);


	not MGM_G98(MGM_W80,E$delay);


	and MGM_G99(MGM_W81,MGM_W80,MGM_W79);


	and MGM_G100(MGM_W82,SD$delay,MGM_W81);


	and MGM_G101(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G102(MGM_W83,D$delay);


	and MGM_G103(MGM_W84,E$delay,MGM_W83);


	and MGM_G104(MGM_W85,SD$delay,MGM_W84);


	and MGM_G105(ENABLE_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G106(MGM_W86,E$delay);


	and MGM_G107(MGM_W87,MGM_W86,D$delay);


	and MGM_G108(MGM_W88,SD$delay,MGM_W87);


	and MGM_G109(ENABLE_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W88);


	and MGM_G110(MGM_W89,E$delay,D$delay);


	not MGM_G111(MGM_W90,SD$delay);


	and MGM_G112(MGM_W91,MGM_W90,MGM_W89);


	not MGM_G113(MGM_W92,SE$delay);


	and MGM_G114(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W92,MGM_W91);


	and MGM_G115(MGM_W93,E$delay,D$delay);


	and MGM_G116(MGM_W94,SD$delay,MGM_W93);


	not MGM_G117(MGM_W95,SE$delay);


	and MGM_G118(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W95,MGM_W94);


	and MGM_G119(MGM_W96,E$delay,D$delay);


	and MGM_G120(MGM_W97,SD$delay,MGM_W96);


	and MGM_G121(ENABLE_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W97);


	not MGM_G122(MGM_W98,CK$delay);


	not MGM_G123(MGM_W99,D$delay);


	and MGM_G124(MGM_W100,MGM_W99,MGM_W98);


	not MGM_G125(MGM_W101,E$delay);


	and MGM_G126(MGM_W102,MGM_W101,MGM_W100);


	not MGM_G127(MGM_W103,SD$delay);


	and MGM_G128(MGM_W104,MGM_W103,MGM_W102);


	not MGM_G129(MGM_W105,SE$delay);


	and MGM_G130(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W105,MGM_W104);


	not MGM_G131(MGM_W106,CK$delay);


	not MGM_G132(MGM_W107,D$delay);


	and MGM_G133(MGM_W108,MGM_W107,MGM_W106);


	not MGM_G134(MGM_W109,E$delay);


	and MGM_G135(MGM_W110,MGM_W109,MGM_W108);


	not MGM_G136(MGM_W111,SD$delay);


	and MGM_G137(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G138(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W112);


	not MGM_G139(MGM_W113,CK$delay);


	not MGM_G140(MGM_W114,D$delay);


	and MGM_G141(MGM_W115,MGM_W114,MGM_W113);


	not MGM_G142(MGM_W116,E$delay);


	and MGM_G143(MGM_W117,MGM_W116,MGM_W115);


	and MGM_G144(MGM_W118,SD$delay,MGM_W117);


	not MGM_G145(MGM_W119,SE$delay);


	and MGM_G146(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W119,MGM_W118);


	not MGM_G147(MGM_W120,CK$delay);


	not MGM_G148(MGM_W121,D$delay);


	and MGM_G149(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G150(MGM_W123,E$delay);


	and MGM_G151(MGM_W124,MGM_W123,MGM_W122);


	and MGM_G152(MGM_W125,SD$delay,MGM_W124);


	and MGM_G153(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W125);


	not MGM_G154(MGM_W126,CK$delay);


	not MGM_G155(MGM_W127,D$delay);


	and MGM_G156(MGM_W128,MGM_W127,MGM_W126);


	and MGM_G157(MGM_W129,E$delay,MGM_W128);


	not MGM_G158(MGM_W130,SD$delay);


	and MGM_G159(MGM_W131,MGM_W130,MGM_W129);


	not MGM_G160(MGM_W132,SE$delay);


	and MGM_G161(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W132,MGM_W131);


	not MGM_G162(MGM_W133,CK$delay);


	not MGM_G163(MGM_W134,D$delay);


	and MGM_G164(MGM_W135,MGM_W134,MGM_W133);


	and MGM_G165(MGM_W136,E$delay,MGM_W135);


	not MGM_G166(MGM_W137,SD$delay);


	and MGM_G167(MGM_W138,MGM_W137,MGM_W136);


	and MGM_G168(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W138);


	not MGM_G169(MGM_W139,CK$delay);


	not MGM_G170(MGM_W140,D$delay);


	and MGM_G171(MGM_W141,MGM_W140,MGM_W139);


	and MGM_G172(MGM_W142,E$delay,MGM_W141);


	and MGM_G173(MGM_W143,SD$delay,MGM_W142);


	not MGM_G174(MGM_W144,SE$delay);


	and MGM_G175(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W144,MGM_W143);


	not MGM_G176(MGM_W145,CK$delay);


	not MGM_G177(MGM_W146,D$delay);


	and MGM_G178(MGM_W147,MGM_W146,MGM_W145);


	and MGM_G179(MGM_W148,E$delay,MGM_W147);


	and MGM_G180(MGM_W149,SD$delay,MGM_W148);


	and MGM_G181(ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W149);


	not MGM_G182(MGM_W150,CK$delay);


	and MGM_G183(MGM_W151,D$delay,MGM_W150);


	not MGM_G184(MGM_W152,E$delay);


	and MGM_G185(MGM_W153,MGM_W152,MGM_W151);


	not MGM_G186(MGM_W154,SD$delay);


	and MGM_G187(MGM_W155,MGM_W154,MGM_W153);


	not MGM_G188(MGM_W156,SE$delay);


	and MGM_G189(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W156,MGM_W155);


	not MGM_G190(MGM_W157,CK$delay);


	and MGM_G191(MGM_W158,D$delay,MGM_W157);


	not MGM_G192(MGM_W159,E$delay);


	and MGM_G193(MGM_W160,MGM_W159,MGM_W158);


	not MGM_G194(MGM_W161,SD$delay);


	and MGM_G195(MGM_W162,MGM_W161,MGM_W160);


	and MGM_G196(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W162);


	not MGM_G197(MGM_W163,CK$delay);


	and MGM_G198(MGM_W164,D$delay,MGM_W163);


	not MGM_G199(MGM_W165,E$delay);


	and MGM_G200(MGM_W166,MGM_W165,MGM_W164);


	and MGM_G201(MGM_W167,SD$delay,MGM_W166);


	not MGM_G202(MGM_W168,SE$delay);


	and MGM_G203(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W168,MGM_W167);


	not MGM_G204(MGM_W169,CK$delay);


	and MGM_G205(MGM_W170,D$delay,MGM_W169);


	not MGM_G206(MGM_W171,E$delay);


	and MGM_G207(MGM_W172,MGM_W171,MGM_W170);


	and MGM_G208(MGM_W173,SD$delay,MGM_W172);


	and MGM_G209(ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W173);


	not MGM_G210(MGM_W174,CK$delay);


	and MGM_G211(MGM_W175,D$delay,MGM_W174);


	and MGM_G212(MGM_W176,E$delay,MGM_W175);


	not MGM_G213(MGM_W177,SD$delay);


	and MGM_G214(MGM_W178,MGM_W177,MGM_W176);


	not MGM_G215(MGM_W179,SE$delay);


	and MGM_G216(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W179,MGM_W178);


	not MGM_G217(MGM_W180,CK$delay);


	and MGM_G218(MGM_W181,D$delay,MGM_W180);


	and MGM_G219(MGM_W182,E$delay,MGM_W181);


	not MGM_G220(MGM_W183,SD$delay);


	and MGM_G221(MGM_W184,MGM_W183,MGM_W182);


	and MGM_G222(ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W184);


	not MGM_G223(MGM_W185,CK$delay);


	and MGM_G224(MGM_W186,D$delay,MGM_W185);


	and MGM_G225(MGM_W187,E$delay,MGM_W186);


	and MGM_G226(MGM_W188,SD$delay,MGM_W187);


	not MGM_G227(MGM_W189,SE$delay);


	and MGM_G228(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W189,MGM_W188);


	not MGM_G229(MGM_W190,CK$delay);


	and MGM_G230(MGM_W191,D$delay,MGM_W190);


	and MGM_G231(MGM_W192,E$delay,MGM_W191);


	and MGM_G232(MGM_W193,SD$delay,MGM_W192);


	and MGM_G233(ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W193);


	not MGM_G234(MGM_W194,D$delay);


	and MGM_G235(MGM_W195,MGM_W194,CK$delay);


	not MGM_G236(MGM_W196,E$delay);


	and MGM_G237(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G238(MGM_W198,SD$delay);


	and MGM_G239(MGM_W199,MGM_W198,MGM_W197);


	not MGM_G240(MGM_W200,SE$delay);


	and MGM_G241(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W200,MGM_W199);


	not MGM_G242(MGM_W201,D$delay);


	and MGM_G243(MGM_W202,MGM_W201,CK$delay);


	not MGM_G244(MGM_W203,E$delay);


	and MGM_G245(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G246(MGM_W205,SD$delay);


	and MGM_G247(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G248(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W206);


	not MGM_G249(MGM_W207,D$delay);


	and MGM_G250(MGM_W208,MGM_W207,CK$delay);


	not MGM_G251(MGM_W209,E$delay);


	and MGM_G252(MGM_W210,MGM_W209,MGM_W208);


	and MGM_G253(MGM_W211,SD$delay,MGM_W210);


	not MGM_G254(MGM_W212,SE$delay);


	and MGM_G255(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W212,MGM_W211);


	not MGM_G256(MGM_W213,D$delay);


	and MGM_G257(MGM_W214,MGM_W213,CK$delay);


	not MGM_G258(MGM_W215,E$delay);


	and MGM_G259(MGM_W216,MGM_W215,MGM_W214);


	and MGM_G260(MGM_W217,SD$delay,MGM_W216);


	and MGM_G261(ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,D$delay);


	and MGM_G263(MGM_W219,MGM_W218,CK$delay);


	and MGM_G264(MGM_W220,E$delay,MGM_W219);


	not MGM_G265(MGM_W221,SD$delay);


	and MGM_G266(MGM_W222,MGM_W221,MGM_W220);


	not MGM_G267(MGM_W223,SE$delay);


	and MGM_G268(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W223,MGM_W222);


	not MGM_G269(MGM_W224,D$delay);


	and MGM_G270(MGM_W225,MGM_W224,CK$delay);


	and MGM_G271(MGM_W226,E$delay,MGM_W225);


	not MGM_G272(MGM_W227,SD$delay);


	and MGM_G273(MGM_W228,MGM_W227,MGM_W226);


	and MGM_G274(ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W228);


	not MGM_G275(MGM_W229,D$delay);


	and MGM_G276(MGM_W230,MGM_W229,CK$delay);


	and MGM_G277(MGM_W231,E$delay,MGM_W230);


	and MGM_G278(MGM_W232,SD$delay,MGM_W231);


	not MGM_G279(MGM_W233,SE$delay);


	and MGM_G280(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G281(MGM_W234,D$delay);


	and MGM_G282(MGM_W235,MGM_W234,CK$delay);


	and MGM_G283(MGM_W236,E$delay,MGM_W235);


	and MGM_G284(MGM_W237,SD$delay,MGM_W236);


	and MGM_G285(ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W237);


	and MGM_G286(MGM_W238,D$delay,CK$delay);


	not MGM_G287(MGM_W239,E$delay);


	and MGM_G288(MGM_W240,MGM_W239,MGM_W238);


	not MGM_G289(MGM_W241,SD$delay);


	and MGM_G290(MGM_W242,MGM_W241,MGM_W240);


	not MGM_G291(MGM_W243,SE$delay);


	and MGM_G292(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W243,MGM_W242);


	and MGM_G293(MGM_W244,D$delay,CK$delay);


	not MGM_G294(MGM_W245,E$delay);


	and MGM_G295(MGM_W246,MGM_W245,MGM_W244);


	not MGM_G296(MGM_W247,SD$delay);


	and MGM_G297(MGM_W248,MGM_W247,MGM_W246);


	and MGM_G298(ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W248);


	and MGM_G299(MGM_W249,D$delay,CK$delay);


	not MGM_G300(MGM_W250,E$delay);


	and MGM_G301(MGM_W251,MGM_W250,MGM_W249);


	and MGM_G302(MGM_W252,SD$delay,MGM_W251);


	not MGM_G303(MGM_W253,SE$delay);


	and MGM_G304(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W253,MGM_W252);


	and MGM_G305(MGM_W254,D$delay,CK$delay);


	not MGM_G306(MGM_W255,E$delay);


	and MGM_G307(MGM_W256,MGM_W255,MGM_W254);


	and MGM_G308(MGM_W257,SD$delay,MGM_W256);


	and MGM_G309(ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE,SE$delay,MGM_W257);


	and MGM_G310(MGM_W258,D$delay,CK$delay);


	and MGM_G311(MGM_W259,E$delay,MGM_W258);


	not MGM_G312(MGM_W260,SD$delay);


	and MGM_G313(MGM_W261,MGM_W260,MGM_W259);


	not MGM_G314(MGM_W262,SE$delay);


	and MGM_G315(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W262,MGM_W261);


	and MGM_G316(MGM_W263,D$delay,CK$delay);


	and MGM_G317(MGM_W264,E$delay,MGM_W263);


	not MGM_G318(MGM_W265,SD$delay);


	and MGM_G319(MGM_W266,MGM_W265,MGM_W264);


	and MGM_G320(ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE,SE$delay,MGM_W266);


	and MGM_G321(MGM_W267,D$delay,CK$delay);


	and MGM_G322(MGM_W268,E$delay,MGM_W267);


	and MGM_G323(MGM_W269,SD$delay,MGM_W268);


	not MGM_G324(MGM_W270,SE$delay);


	and MGM_G325(ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE,MGM_W270,MGM_W269);


	and MGM_G326(MGM_W271,D$delay,CK$delay);


	and MGM_G327(MGM_W272,E$delay,MGM_W271);


	and MGM_G328(MGM_W273,SD$delay,MGM_W272);


	and MGM_G329(ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE,SE$delay,MGM_W273);


	not MGM_G330(MGM_W274,D$delay);


	not MGM_G331(MGM_W275,E$delay);


	and MGM_G332(MGM_W276,MGM_W275,MGM_W274);


	and MGM_G333(MGM_W277,RB$delay,MGM_W276);


	and MGM_G334(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W277);


	not MGM_G335(MGM_W278,D$delay);


	and MGM_G336(MGM_W279,E$delay,MGM_W278);


	and MGM_G337(MGM_W280,RB$delay,MGM_W279);


	and MGM_G338(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W280);


	not MGM_G339(MGM_W281,E$delay);


	and MGM_G340(MGM_W282,MGM_W281,D$delay);


	and MGM_G341(MGM_W283,RB$delay,MGM_W282);


	and MGM_G342(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W283);


	and MGM_G343(MGM_W284,E$delay,D$delay);


	and MGM_G344(MGM_W285,RB$delay,MGM_W284);


	and MGM_G345(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W285);


	not MGM_G346(MGM_W286,D$delay);


	not MGM_G347(MGM_W287,E$delay);


	and MGM_G348(MGM_W288,MGM_W287,MGM_W286);


	and MGM_G349(MGM_W289,RB$delay,MGM_W288);


	not MGM_G350(MGM_W290,SD$delay);


	and MGM_G351(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W290,MGM_W289);


	not MGM_G352(MGM_W291,D$delay);


	not MGM_G353(MGM_W292,E$delay);


	and MGM_G354(MGM_W293,MGM_W292,MGM_W291);


	and MGM_G355(MGM_W294,RB$delay,MGM_W293);


	and MGM_G356(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W294);


	not MGM_G357(MGM_W295,D$delay);


	and MGM_G358(MGM_W296,E$delay,MGM_W295);


	and MGM_G359(MGM_W297,RB$delay,MGM_W296);


	and MGM_G360(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W297);


	not MGM_G361(MGM_W298,E$delay);


	and MGM_G362(MGM_W299,MGM_W298,D$delay);


	and MGM_G363(MGM_W300,RB$delay,MGM_W299);


	not MGM_G364(MGM_W301,SD$delay);


	and MGM_G365(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W301,MGM_W300);


	not MGM_G366(MGM_W302,E$delay);


	and MGM_G367(MGM_W303,MGM_W302,D$delay);


	and MGM_G368(MGM_W304,RB$delay,MGM_W303);


	and MGM_G369(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W304);


	and MGM_G370(MGM_W305,E$delay,D$delay);


	and MGM_G371(MGM_W306,RB$delay,MGM_W305);


	not MGM_G372(MGM_W307,SD$delay);


	and MGM_G373(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W307,MGM_W306);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_E_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEZRM1HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM1HM_func SDFEZRM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEZRM1HM_func SDFEZRM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEZRM2HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM2HM_func SDFEZRM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEZRM2HM_func SDFEZRM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEZRM4HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM4HM_func SDFEZRM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEZRM4HM_func SDFEZRM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFEZRM8HM( Q, QB, CK, D, E, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM8HM_func SDFEZRM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.E(E),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire E$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFEZRM8HM_func SDFEZRM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.E(E$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,E$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,RB$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D$delay);


	not MGM_G10(MGM_W9,E$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,RB$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D$delay);


	not MGM_G18(MGM_W16,E$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,RB$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D$delay);


	not MGM_G26(MGM_W23,E$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,RB$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D$delay);


	not MGM_G33(MGM_W29,E$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,RB$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	and MGM_G38(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W33);


	not MGM_G39(MGM_W34,D$delay);


	not MGM_G40(MGM_W35,E$delay);


	and MGM_G41(MGM_W36,MGM_W35,MGM_W34);


	and MGM_G42(MGM_W37,RB$delay,MGM_W36);


	and MGM_G43(MGM_W38,SD$delay,MGM_W37);


	and MGM_G44(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W38);


	not MGM_G45(MGM_W39,D$delay);


	and MGM_G46(MGM_W40,E$delay,MGM_W39);


	not MGM_G47(MGM_W41,RB$delay);


	and MGM_G48(MGM_W42,MGM_W41,MGM_W40);


	not MGM_G49(MGM_W43,SD$delay);


	and MGM_G50(MGM_W44,MGM_W43,MGM_W42);


	not MGM_G51(MGM_W45,SE$delay);


	and MGM_G52(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W45,MGM_W44);


	not MGM_G53(MGM_W46,D$delay);


	and MGM_G54(MGM_W47,E$delay,MGM_W46);


	not MGM_G55(MGM_W48,RB$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G57(MGM_W50,SD$delay);


	and MGM_G58(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G59(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D$delay);


	and MGM_G61(MGM_W53,E$delay,MGM_W52);


	not MGM_G62(MGM_W54,RB$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G64(MGM_W56,SD$delay,MGM_W55);


	not MGM_G65(MGM_W57,SE$delay);


	and MGM_G66(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W57,MGM_W56);


	not MGM_G67(MGM_W58,D$delay);


	and MGM_G68(MGM_W59,E$delay,MGM_W58);


	not MGM_G69(MGM_W60,RB$delay);


	and MGM_G70(MGM_W61,MGM_W60,MGM_W59);


	and MGM_G71(MGM_W62,SD$delay,MGM_W61);


	and MGM_G72(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W62);


	not MGM_G73(MGM_W63,D$delay);


	and MGM_G74(MGM_W64,E$delay,MGM_W63);


	and MGM_G75(MGM_W65,RB$delay,MGM_W64);


	not MGM_G76(MGM_W66,SD$delay);


	and MGM_G77(MGM_W67,MGM_W66,MGM_W65);


	not MGM_G78(MGM_W68,SE$delay);


	and MGM_G79(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G80(MGM_W69,D$delay);


	and MGM_G81(MGM_W70,E$delay,MGM_W69);


	and MGM_G82(MGM_W71,RB$delay,MGM_W70);


	not MGM_G83(MGM_W72,SD$delay);


	and MGM_G84(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G85(ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G86(MGM_W74,D$delay);


	and MGM_G87(MGM_W75,E$delay,MGM_W74);


	and MGM_G88(MGM_W76,RB$delay,MGM_W75);


	and MGM_G89(MGM_W77,SD$delay,MGM_W76);


	not MGM_G90(MGM_W78,SE$delay);


	and MGM_G91(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W78,MGM_W77);


	not MGM_G92(MGM_W79,D$delay);


	and MGM_G93(MGM_W80,E$delay,MGM_W79);


	and MGM_G94(MGM_W81,RB$delay,MGM_W80);


	and MGM_G95(MGM_W82,SD$delay,MGM_W81);


	and MGM_G96(ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W82);


	not MGM_G97(MGM_W83,E$delay);


	and MGM_G98(MGM_W84,MGM_W83,D$delay);


	not MGM_G99(MGM_W85,RB$delay);


	and MGM_G100(MGM_W86,MGM_W85,MGM_W84);


	not MGM_G101(MGM_W87,SD$delay);


	and MGM_G102(MGM_W88,MGM_W87,MGM_W86);


	not MGM_G103(MGM_W89,SE$delay);


	and MGM_G104(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G105(MGM_W90,E$delay);


	and MGM_G106(MGM_W91,MGM_W90,D$delay);


	not MGM_G107(MGM_W92,RB$delay);


	and MGM_G108(MGM_W93,MGM_W92,MGM_W91);


	not MGM_G109(MGM_W94,SD$delay);


	and MGM_G110(MGM_W95,MGM_W94,MGM_W93);


	and MGM_G111(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,E$delay);


	and MGM_G113(MGM_W97,MGM_W96,D$delay);


	not MGM_G114(MGM_W98,RB$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G116(MGM_W100,SD$delay,MGM_W99);


	not MGM_G117(MGM_W101,SE$delay);


	and MGM_G118(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W101,MGM_W100);


	not MGM_G119(MGM_W102,E$delay);


	and MGM_G120(MGM_W103,MGM_W102,D$delay);


	not MGM_G121(MGM_W104,RB$delay);


	and MGM_G122(MGM_W105,MGM_W104,MGM_W103);


	and MGM_G123(MGM_W106,SD$delay,MGM_W105);


	and MGM_G124(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W106);


	not MGM_G125(MGM_W107,E$delay);


	and MGM_G126(MGM_W108,MGM_W107,D$delay);


	and MGM_G127(MGM_W109,RB$delay,MGM_W108);


	not MGM_G128(MGM_W110,SD$delay);


	and MGM_G129(MGM_W111,MGM_W110,MGM_W109);


	and MGM_G130(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W111);


	not MGM_G131(MGM_W112,E$delay);


	and MGM_G132(MGM_W113,MGM_W112,D$delay);


	and MGM_G133(MGM_W114,RB$delay,MGM_W113);


	and MGM_G134(MGM_W115,SD$delay,MGM_W114);


	and MGM_G135(ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W115);


	and MGM_G136(MGM_W116,E$delay,D$delay);


	not MGM_G137(MGM_W117,RB$delay);


	and MGM_G138(MGM_W118,MGM_W117,MGM_W116);


	not MGM_G139(MGM_W119,SD$delay);


	and MGM_G140(MGM_W120,MGM_W119,MGM_W118);


	not MGM_G141(MGM_W121,SE$delay);


	and MGM_G142(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W121,MGM_W120);


	and MGM_G143(MGM_W122,E$delay,D$delay);


	not MGM_G144(MGM_W123,RB$delay);


	and MGM_G145(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G146(MGM_W125,SD$delay);


	and MGM_G147(MGM_W126,MGM_W125,MGM_W124);


	and MGM_G148(ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W126);


	and MGM_G149(MGM_W127,E$delay,D$delay);


	not MGM_G150(MGM_W128,RB$delay);


	and MGM_G151(MGM_W129,MGM_W128,MGM_W127);


	and MGM_G152(MGM_W130,SD$delay,MGM_W129);


	not MGM_G153(MGM_W131,SE$delay);


	and MGM_G154(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G155(MGM_W132,E$delay,D$delay);


	not MGM_G156(MGM_W133,RB$delay);


	and MGM_G157(MGM_W134,MGM_W133,MGM_W132);


	and MGM_G158(MGM_W135,SD$delay,MGM_W134);


	and MGM_G159(ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W135);


	and MGM_G160(MGM_W136,E$delay,D$delay);


	and MGM_G161(MGM_W137,RB$delay,MGM_W136);


	not MGM_G162(MGM_W138,SD$delay);


	and MGM_G163(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G164(MGM_W140,SE$delay);


	and MGM_G165(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	and MGM_G166(MGM_W141,E$delay,D$delay);


	and MGM_G167(MGM_W142,RB$delay,MGM_W141);


	not MGM_G168(MGM_W143,SD$delay);


	and MGM_G169(MGM_W144,MGM_W143,MGM_W142);


	and MGM_G170(ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W144);


	and MGM_G171(MGM_W145,E$delay,D$delay);


	and MGM_G172(MGM_W146,RB$delay,MGM_W145);


	and MGM_G173(MGM_W147,SD$delay,MGM_W146);


	not MGM_G174(MGM_W148,SE$delay);


	and MGM_G175(ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W148,MGM_W147);


	and MGM_G176(MGM_W149,E$delay,D$delay);


	and MGM_G177(MGM_W150,RB$delay,MGM_W149);


	and MGM_G178(MGM_W151,SD$delay,MGM_W150);


	and MGM_G179(ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W151);


	and MGM_G180(MGM_W152,RB$delay,E$delay);


	not MGM_G181(MGM_W153,SD$delay);


	and MGM_G182(MGM_W154,MGM_W153,MGM_W152);


	not MGM_G183(MGM_W155,SE$delay);


	and MGM_G184(ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G185(MGM_W156,RB$delay,E$delay);


	and MGM_G186(MGM_W157,SD$delay,MGM_W156);


	not MGM_G187(MGM_W158,SE$delay);


	and MGM_G188(ENABLE_E_AND_RB_AND_SD_AND_NOT_SE,MGM_W158,MGM_W157);


	not MGM_G189(MGM_W159,D$delay);


	and MGM_G190(MGM_W160,RB$delay,MGM_W159);


	not MGM_G191(MGM_W161,SD$delay);


	and MGM_G192(MGM_W162,MGM_W161,MGM_W160);


	not MGM_G193(MGM_W163,SE$delay);


	and MGM_G194(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W163,MGM_W162);


	not MGM_G195(MGM_W164,D$delay);


	and MGM_G196(MGM_W165,RB$delay,MGM_W164);


	and MGM_G197(MGM_W166,SD$delay,MGM_W165);


	not MGM_G198(MGM_W167,SE$delay);


	and MGM_G199(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	and MGM_G200(MGM_W168,RB$delay,D$delay);


	not MGM_G201(MGM_W169,SD$delay);


	and MGM_G202(MGM_W170,MGM_W169,MGM_W168);


	not MGM_G203(MGM_W171,SE$delay);


	and MGM_G204(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W171,MGM_W170);


	and MGM_G205(MGM_W172,RB$delay,D$delay);


	and MGM_G206(MGM_W173,SD$delay,MGM_W172);


	not MGM_G207(MGM_W174,SE$delay);


	and MGM_G208(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W174,MGM_W173);


	not MGM_G209(MGM_W175,D$delay);


	not MGM_G210(MGM_W176,E$delay);


	and MGM_G211(MGM_W177,MGM_W176,MGM_W175);


	not MGM_G212(MGM_W178,SD$delay);


	and MGM_G213(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G214(MGM_W180,SE$delay);


	and MGM_G215(ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G216(MGM_W181,D$delay);


	not MGM_G217(MGM_W182,E$delay);


	and MGM_G218(MGM_W183,MGM_W182,MGM_W181);


	and MGM_G219(MGM_W184,SD$delay,MGM_W183);


	not MGM_G220(MGM_W185,SE$delay);


	and MGM_G221(ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W185,MGM_W184);


	not MGM_G222(MGM_W186,E$delay);


	and MGM_G223(MGM_W187,MGM_W186,D$delay);


	not MGM_G224(MGM_W188,SD$delay);


	and MGM_G225(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G226(MGM_W190,SE$delay);


	and MGM_G227(ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	not MGM_G228(MGM_W191,E$delay);


	and MGM_G229(MGM_W192,MGM_W191,D$delay);


	and MGM_G230(MGM_W193,SD$delay,MGM_W192);


	not MGM_G231(MGM_W194,SE$delay);


	and MGM_G232(ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE,MGM_W194,MGM_W193);


	and MGM_G233(MGM_W195,E$delay,D$delay);


	not MGM_G234(MGM_W196,SD$delay);


	and MGM_G235(MGM_W197,MGM_W196,MGM_W195);


	not MGM_G236(MGM_W198,SE$delay);


	and MGM_G237(ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE,MGM_W198,MGM_W197);


	and MGM_G238(MGM_W199,E$delay,D$delay);


	and MGM_G239(MGM_W200,SD$delay,MGM_W199);


	not MGM_G240(MGM_W201,SE$delay);


	and MGM_G241(ENABLE_D_AND_E_AND_SD_AND_NOT_SE,MGM_W201,MGM_W200);


	not MGM_G242(MGM_W202,D$delay);


	not MGM_G243(MGM_W203,E$delay);


	and MGM_G244(MGM_W204,MGM_W203,MGM_W202);


	not MGM_G245(MGM_W205,RB$delay);


	and MGM_G246(MGM_W206,MGM_W205,MGM_W204);


	and MGM_G247(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W206);


	not MGM_G248(MGM_W207,D$delay);


	not MGM_G249(MGM_W208,E$delay);


	and MGM_G250(MGM_W209,MGM_W208,MGM_W207);


	and MGM_G251(MGM_W210,RB$delay,MGM_W209);


	and MGM_G252(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W210);


	not MGM_G253(MGM_W211,D$delay);


	and MGM_G254(MGM_W212,E$delay,MGM_W211);


	not MGM_G255(MGM_W213,RB$delay);


	and MGM_G256(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G257(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W214);


	not MGM_G258(MGM_W215,D$delay);


	and MGM_G259(MGM_W216,E$delay,MGM_W215);


	and MGM_G260(MGM_W217,RB$delay,MGM_W216);


	and MGM_G261(ENABLE_NOT_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W217);


	not MGM_G262(MGM_W218,E$delay);


	and MGM_G263(MGM_W219,MGM_W218,D$delay);


	not MGM_G264(MGM_W220,RB$delay);


	and MGM_G265(MGM_W221,MGM_W220,MGM_W219);


	and MGM_G266(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W221);


	not MGM_G267(MGM_W222,E$delay);


	and MGM_G268(MGM_W223,MGM_W222,D$delay);


	and MGM_G269(MGM_W224,RB$delay,MGM_W223);


	and MGM_G270(ENABLE_D_AND_NOT_E_AND_RB_AND_SE,SE$delay,MGM_W224);


	and MGM_G271(MGM_W225,E$delay,D$delay);


	not MGM_G272(MGM_W226,RB$delay);


	and MGM_G273(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G274(ENABLE_D_AND_E_AND_NOT_RB_AND_SE,SE$delay,MGM_W227);


	and MGM_G275(MGM_W228,E$delay,D$delay);


	and MGM_G276(MGM_W229,RB$delay,MGM_W228);


	and MGM_G277(ENABLE_D_AND_E_AND_RB_AND_SE,SE$delay,MGM_W229);


	not MGM_G278(MGM_W230,D$delay);


	not MGM_G279(MGM_W231,E$delay);


	and MGM_G280(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G281(MGM_W233,RB$delay);


	and MGM_G282(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G283(ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W234);


	not MGM_G284(MGM_W235,D$delay);


	not MGM_G285(MGM_W236,E$delay);


	and MGM_G286(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G287(MGM_W238,RB$delay,MGM_W237);


	not MGM_G288(MGM_W239,SD$delay);


	and MGM_G289(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W239,MGM_W238);


	not MGM_G290(MGM_W240,D$delay);


	not MGM_G291(MGM_W241,E$delay);


	and MGM_G292(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G293(MGM_W243,RB$delay,MGM_W242);


	and MGM_G294(ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W243);


	not MGM_G295(MGM_W244,D$delay);


	and MGM_G296(MGM_W245,E$delay,MGM_W244);


	not MGM_G297(MGM_W246,RB$delay);


	and MGM_G298(MGM_W247,MGM_W246,MGM_W245);


	and MGM_G299(ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W247);


	not MGM_G300(MGM_W248,D$delay);


	and MGM_G301(MGM_W249,E$delay,MGM_W248);


	and MGM_G302(MGM_W250,RB$delay,MGM_W249);


	and MGM_G303(ENABLE_NOT_D_AND_E_AND_RB_AND_SD,SD$delay,MGM_W250);


	not MGM_G304(MGM_W251,E$delay);


	and MGM_G305(MGM_W252,MGM_W251,D$delay);


	not MGM_G306(MGM_W253,RB$delay);


	and MGM_G307(MGM_W254,MGM_W253,MGM_W252);


	and MGM_G308(ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W254);


	not MGM_G309(MGM_W255,E$delay);


	and MGM_G310(MGM_W256,MGM_W255,D$delay);


	and MGM_G311(MGM_W257,RB$delay,MGM_W256);


	not MGM_G312(MGM_W258,SD$delay);


	and MGM_G313(ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD,MGM_W258,MGM_W257);


	not MGM_G314(MGM_W259,E$delay);


	and MGM_G315(MGM_W260,MGM_W259,D$delay);


	and MGM_G316(MGM_W261,RB$delay,MGM_W260);


	and MGM_G317(ENABLE_D_AND_NOT_E_AND_RB_AND_SD,SD$delay,MGM_W261);


	and MGM_G318(MGM_W262,E$delay,D$delay);


	not MGM_G319(MGM_W263,RB$delay);


	and MGM_G320(MGM_W264,MGM_W263,MGM_W262);


	and MGM_G321(ENABLE_D_AND_E_AND_NOT_RB_AND_SD,SD$delay,MGM_W264);


	and MGM_G322(MGM_W265,E$delay,D$delay);


	and MGM_G323(MGM_W266,RB$delay,MGM_W265);


	not MGM_G324(MGM_W267,SD$delay);


	and MGM_G325(ENABLE_D_AND_E_AND_RB_AND_NOT_SD,MGM_W267,MGM_W266);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_E_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_E_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_E_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_E_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFM1HM( Q, QB, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFM1HM_func SDFM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFM1HM_func SDFM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFM2HM( Q, QB, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFM2HM_func SDFM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFM2HM_func SDFM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFM4HM( Q, QB, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFM4HM_func SDFM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFM4HM_func SDFM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFM8HM( Q, QB, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFM8HM_func SDFM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFM8HM_func SDFM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMM1HM( Q, QB, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMM1HM_func SDFMM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMM1HM_func SDFMM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMM2HM( Q, QB, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMM2HM_func SDFMM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMM2HM_func SDFMM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMM4HM( Q, QB, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMM4HM_func SDFMM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMM4HM_func SDFMM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMM8HM( Q, QB, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMM8HM_func SDFMM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMM8HM_func SDFMM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMQM1HM( Q, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMQM1HM_func SDFMQM1HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMQM1HM_func SDFMQM1HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMQM2HM( Q, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMQM2HM_func SDFMQM2HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMQM2HM_func SDFMQM2HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMQM4HM( Q, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMQM4HM_func SDFMQM4HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMQM4HM_func SDFMQM4HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFMQM8HM( Q, CK, D1, D2, S, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFMQM8HM_func SDFMQM8HM_behav_inst(.Q(Q),.CK(CK),.D1(D1),.D2(D2),.S(S),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D1$delay ;

	wire D2$delay ;

	wire S$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFMQM8HM_func SDFMQM8HM_inst(.Q(Q),.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D1$delay);


	not MGM_G1(MGM_W1,D2$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,S$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SD$delay);


	and MGM_G6(MGM_W6,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W7,SE$delay);


	and MGM_G8(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W7,MGM_W6);


	not MGM_G9(MGM_W8,D1$delay);


	not MGM_G10(MGM_W9,D2$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	not MGM_G12(MGM_W11,S$delay);


	and MGM_G13(MGM_W12,MGM_W11,MGM_W10);


	not MGM_G14(MGM_W13,SD$delay);


	and MGM_G15(MGM_W14,MGM_W13,MGM_W12);


	and MGM_G16(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W14);


	not MGM_G17(MGM_W15,D1$delay);


	not MGM_G18(MGM_W16,D2$delay);


	and MGM_G19(MGM_W17,MGM_W16,MGM_W15);


	not MGM_G20(MGM_W18,S$delay);


	and MGM_G21(MGM_W19,MGM_W18,MGM_W17);


	and MGM_G22(MGM_W20,SD$delay,MGM_W19);


	not MGM_G23(MGM_W21,SE$delay);


	and MGM_G24(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G25(MGM_W22,D1$delay);


	not MGM_G26(MGM_W23,D2$delay);


	and MGM_G27(MGM_W24,MGM_W23,MGM_W22);


	not MGM_G28(MGM_W25,S$delay);


	and MGM_G29(MGM_W26,MGM_W25,MGM_W24);


	and MGM_G30(MGM_W27,SD$delay,MGM_W26);


	and MGM_G31(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G32(MGM_W28,D1$delay);


	not MGM_G33(MGM_W29,D2$delay);


	and MGM_G34(MGM_W30,MGM_W29,MGM_W28);


	and MGM_G35(MGM_W31,S$delay,MGM_W30);


	not MGM_G36(MGM_W32,SD$delay);


	and MGM_G37(MGM_W33,MGM_W32,MGM_W31);


	not MGM_G38(MGM_W34,SE$delay);


	and MGM_G39(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W34,MGM_W33);


	not MGM_G40(MGM_W35,D1$delay);


	not MGM_G41(MGM_W36,D2$delay);


	and MGM_G42(MGM_W37,MGM_W36,MGM_W35);


	and MGM_G43(MGM_W38,S$delay,MGM_W37);


	not MGM_G44(MGM_W39,SD$delay);


	and MGM_G45(MGM_W40,MGM_W39,MGM_W38);


	and MGM_G46(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G47(MGM_W41,D1$delay);


	not MGM_G48(MGM_W42,D2$delay);


	and MGM_G49(MGM_W43,MGM_W42,MGM_W41);


	and MGM_G50(MGM_W44,S$delay,MGM_W43);


	and MGM_G51(MGM_W45,SD$delay,MGM_W44);


	not MGM_G52(MGM_W46,SE$delay);


	and MGM_G53(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G54(MGM_W47,D1$delay);


	not MGM_G55(MGM_W48,D2$delay);


	and MGM_G56(MGM_W49,MGM_W48,MGM_W47);


	and MGM_G57(MGM_W50,S$delay,MGM_W49);


	and MGM_G58(MGM_W51,SD$delay,MGM_W50);


	and MGM_G59(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G60(MGM_W52,D1$delay);


	and MGM_G61(MGM_W53,D2$delay,MGM_W52);


	not MGM_G62(MGM_W54,S$delay);


	and MGM_G63(MGM_W55,MGM_W54,MGM_W53);


	not MGM_G64(MGM_W56,SD$delay);


	and MGM_G65(MGM_W57,MGM_W56,MGM_W55);


	not MGM_G66(MGM_W58,SE$delay);


	and MGM_G67(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W58,MGM_W57);


	not MGM_G68(MGM_W59,D1$delay);


	and MGM_G69(MGM_W60,D2$delay,MGM_W59);


	not MGM_G70(MGM_W61,S$delay);


	and MGM_G71(MGM_W62,MGM_W61,MGM_W60);


	not MGM_G72(MGM_W63,SD$delay);


	and MGM_G73(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G74(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G75(MGM_W65,D1$delay);


	and MGM_G76(MGM_W66,D2$delay,MGM_W65);


	not MGM_G77(MGM_W67,S$delay);


	and MGM_G78(MGM_W68,MGM_W67,MGM_W66);


	and MGM_G79(MGM_W69,SD$delay,MGM_W68);


	not MGM_G80(MGM_W70,SE$delay);


	and MGM_G81(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W70,MGM_W69);


	not MGM_G82(MGM_W71,D1$delay);


	and MGM_G83(MGM_W72,D2$delay,MGM_W71);


	not MGM_G84(MGM_W73,S$delay);


	and MGM_G85(MGM_W74,MGM_W73,MGM_W72);


	and MGM_G86(MGM_W75,SD$delay,MGM_W74);


	and MGM_G87(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W75);


	not MGM_G88(MGM_W76,D1$delay);


	and MGM_G89(MGM_W77,D2$delay,MGM_W76);


	and MGM_G90(MGM_W78,S$delay,MGM_W77);


	not MGM_G91(MGM_W79,SD$delay);


	and MGM_G92(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G93(MGM_W81,SE$delay);


	and MGM_G94(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G95(MGM_W82,D1$delay);


	and MGM_G96(MGM_W83,D2$delay,MGM_W82);


	and MGM_G97(MGM_W84,S$delay,MGM_W83);


	not MGM_G98(MGM_W85,SD$delay);


	and MGM_G99(MGM_W86,MGM_W85,MGM_W84);


	and MGM_G100(ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W86);


	not MGM_G101(MGM_W87,D1$delay);


	and MGM_G102(MGM_W88,D2$delay,MGM_W87);


	and MGM_G103(MGM_W89,S$delay,MGM_W88);


	and MGM_G104(MGM_W90,SD$delay,MGM_W89);


	not MGM_G105(MGM_W91,SE$delay);


	and MGM_G106(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W91,MGM_W90);


	not MGM_G107(MGM_W92,D1$delay);


	and MGM_G108(MGM_W93,D2$delay,MGM_W92);


	and MGM_G109(MGM_W94,S$delay,MGM_W93);


	and MGM_G110(MGM_W95,SD$delay,MGM_W94);


	and MGM_G111(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W95);


	not MGM_G112(MGM_W96,D2$delay);


	and MGM_G113(MGM_W97,MGM_W96,D1$delay);


	not MGM_G114(MGM_W98,S$delay);


	and MGM_G115(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G116(MGM_W100,SD$delay);


	and MGM_G117(MGM_W101,MGM_W100,MGM_W99);


	not MGM_G118(MGM_W102,SE$delay);


	and MGM_G119(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	not MGM_G120(MGM_W103,D2$delay);


	and MGM_G121(MGM_W104,MGM_W103,D1$delay);


	not MGM_G122(MGM_W105,S$delay);


	and MGM_G123(MGM_W106,MGM_W105,MGM_W104);


	not MGM_G124(MGM_W107,SD$delay);


	and MGM_G125(MGM_W108,MGM_W107,MGM_W106);


	and MGM_G126(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G127(MGM_W109,D2$delay);


	and MGM_G128(MGM_W110,MGM_W109,D1$delay);


	not MGM_G129(MGM_W111,S$delay);


	and MGM_G130(MGM_W112,MGM_W111,MGM_W110);


	and MGM_G131(MGM_W113,SD$delay,MGM_W112);


	not MGM_G132(MGM_W114,SE$delay);


	and MGM_G133(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G134(MGM_W115,D2$delay);


	and MGM_G135(MGM_W116,MGM_W115,D1$delay);


	not MGM_G136(MGM_W117,S$delay);


	and MGM_G137(MGM_W118,MGM_W117,MGM_W116);


	and MGM_G138(MGM_W119,SD$delay,MGM_W118);


	and MGM_G139(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W119);


	not MGM_G140(MGM_W120,D2$delay);


	and MGM_G141(MGM_W121,MGM_W120,D1$delay);


	and MGM_G142(MGM_W122,S$delay,MGM_W121);


	not MGM_G143(MGM_W123,SD$delay);


	and MGM_G144(MGM_W124,MGM_W123,MGM_W122);


	not MGM_G145(MGM_W125,SE$delay);


	and MGM_G146(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W125,MGM_W124);


	not MGM_G147(MGM_W126,D2$delay);


	and MGM_G148(MGM_W127,MGM_W126,D1$delay);


	and MGM_G149(MGM_W128,S$delay,MGM_W127);


	not MGM_G150(MGM_W129,SD$delay);


	and MGM_G151(MGM_W130,MGM_W129,MGM_W128);


	and MGM_G152(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W130);


	not MGM_G153(MGM_W131,D2$delay);


	and MGM_G154(MGM_W132,MGM_W131,D1$delay);


	and MGM_G155(MGM_W133,S$delay,MGM_W132);


	and MGM_G156(MGM_W134,SD$delay,MGM_W133);


	not MGM_G157(MGM_W135,SE$delay);


	and MGM_G158(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W135,MGM_W134);


	not MGM_G159(MGM_W136,D2$delay);


	and MGM_G160(MGM_W137,MGM_W136,D1$delay);


	and MGM_G161(MGM_W138,S$delay,MGM_W137);


	and MGM_G162(MGM_W139,SD$delay,MGM_W138);


	and MGM_G163(ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W139);


	and MGM_G164(MGM_W140,D2$delay,D1$delay);


	not MGM_G165(MGM_W141,S$delay);


	and MGM_G166(MGM_W142,MGM_W141,MGM_W140);


	not MGM_G167(MGM_W143,SD$delay);


	and MGM_G168(MGM_W144,MGM_W143,MGM_W142);


	not MGM_G169(MGM_W145,SE$delay);


	and MGM_G170(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W145,MGM_W144);


	and MGM_G171(MGM_W146,D2$delay,D1$delay);


	not MGM_G172(MGM_W147,S$delay);


	and MGM_G173(MGM_W148,MGM_W147,MGM_W146);


	not MGM_G174(MGM_W149,SD$delay);


	and MGM_G175(MGM_W150,MGM_W149,MGM_W148);


	and MGM_G176(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W150);


	and MGM_G177(MGM_W151,D2$delay,D1$delay);


	not MGM_G178(MGM_W152,S$delay);


	and MGM_G179(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G180(MGM_W154,SD$delay,MGM_W153);


	not MGM_G181(MGM_W155,SE$delay);


	and MGM_G182(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W155,MGM_W154);


	and MGM_G183(MGM_W156,D2$delay,D1$delay);


	not MGM_G184(MGM_W157,S$delay);


	and MGM_G185(MGM_W158,MGM_W157,MGM_W156);


	and MGM_G186(MGM_W159,SD$delay,MGM_W158);


	and MGM_G187(ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE,SE$delay,MGM_W159);


	and MGM_G188(MGM_W160,D2$delay,D1$delay);


	and MGM_G189(MGM_W161,S$delay,MGM_W160);


	not MGM_G190(MGM_W162,SD$delay);


	and MGM_G191(MGM_W163,MGM_W162,MGM_W161);


	not MGM_G192(MGM_W164,SE$delay);


	and MGM_G193(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W164,MGM_W163);


	and MGM_G194(MGM_W165,D2$delay,D1$delay);


	and MGM_G195(MGM_W166,S$delay,MGM_W165);


	not MGM_G196(MGM_W167,SD$delay);


	and MGM_G197(MGM_W168,MGM_W167,MGM_W166);


	and MGM_G198(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE,SE$delay,MGM_W168);


	and MGM_G199(MGM_W169,D2$delay,D1$delay);


	and MGM_G200(MGM_W170,S$delay,MGM_W169);


	and MGM_G201(MGM_W171,SD$delay,MGM_W170);


	not MGM_G202(MGM_W172,SE$delay);


	and MGM_G203(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W172,MGM_W171);


	and MGM_G204(MGM_W173,D2$delay,D1$delay);


	and MGM_G205(MGM_W174,S$delay,MGM_W173);


	and MGM_G206(MGM_W175,SD$delay,MGM_W174);


	and MGM_G207(ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE,SE$delay,MGM_W175);


	not MGM_G208(MGM_W176,D2$delay);


	and MGM_G209(MGM_W177,S$delay,MGM_W176);


	not MGM_G210(MGM_W178,SD$delay);


	and MGM_G211(MGM_W179,MGM_W178,MGM_W177);


	not MGM_G212(MGM_W180,SE$delay);


	and MGM_G213(ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W180,MGM_W179);


	not MGM_G214(MGM_W181,D2$delay);


	and MGM_G215(MGM_W182,S$delay,MGM_W181);


	and MGM_G216(MGM_W183,SD$delay,MGM_W182);


	not MGM_G217(MGM_W184,SE$delay);


	and MGM_G218(ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W184,MGM_W183);


	and MGM_G219(MGM_W185,S$delay,D2$delay);


	not MGM_G220(MGM_W186,SD$delay);


	and MGM_G221(MGM_W187,MGM_W186,MGM_W185);


	not MGM_G222(MGM_W188,SE$delay);


	and MGM_G223(ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE,MGM_W188,MGM_W187);


	and MGM_G224(MGM_W189,S$delay,D2$delay);


	and MGM_G225(MGM_W190,SD$delay,MGM_W189);


	not MGM_G226(MGM_W191,SE$delay);


	and MGM_G227(ENABLE_D2_AND_S_AND_SD_AND_NOT_SE,MGM_W191,MGM_W190);


	not MGM_G228(MGM_W192,D1$delay);


	not MGM_G229(MGM_W193,S$delay);


	and MGM_G230(MGM_W194,MGM_W193,MGM_W192);


	not MGM_G231(MGM_W195,SD$delay);


	and MGM_G232(MGM_W196,MGM_W195,MGM_W194);


	not MGM_G233(MGM_W197,SE$delay);


	and MGM_G234(ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W197,MGM_W196);


	not MGM_G235(MGM_W198,D1$delay);


	not MGM_G236(MGM_W199,S$delay);


	and MGM_G237(MGM_W200,MGM_W199,MGM_W198);


	and MGM_G238(MGM_W201,SD$delay,MGM_W200);


	not MGM_G239(MGM_W202,SE$delay);


	and MGM_G240(ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W202,MGM_W201);


	not MGM_G241(MGM_W203,S$delay);


	and MGM_G242(MGM_W204,MGM_W203,D1$delay);


	not MGM_G243(MGM_W205,SD$delay);


	and MGM_G244(MGM_W206,MGM_W205,MGM_W204);


	not MGM_G245(MGM_W207,SE$delay);


	and MGM_G246(ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE,MGM_W207,MGM_W206);


	not MGM_G247(MGM_W208,S$delay);


	and MGM_G248(MGM_W209,MGM_W208,D1$delay);


	and MGM_G249(MGM_W210,SD$delay,MGM_W209);


	not MGM_G250(MGM_W211,SE$delay);


	and MGM_G251(ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	not MGM_G252(MGM_W212,D1$delay);


	and MGM_G253(MGM_W213,D2$delay,MGM_W212);


	not MGM_G254(MGM_W214,SD$delay);


	and MGM_G255(MGM_W215,MGM_W214,MGM_W213);


	not MGM_G256(MGM_W216,SE$delay);


	and MGM_G257(ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE,MGM_W216,MGM_W215);


	not MGM_G258(MGM_W217,D1$delay);


	and MGM_G259(MGM_W218,D2$delay,MGM_W217);


	and MGM_G260(MGM_W219,SD$delay,MGM_W218);


	not MGM_G261(MGM_W220,SE$delay);


	and MGM_G262(ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE,MGM_W220,MGM_W219);


	not MGM_G263(MGM_W221,D2$delay);


	and MGM_G264(MGM_W222,MGM_W221,D1$delay);


	not MGM_G265(MGM_W223,SD$delay);


	and MGM_G266(MGM_W224,MGM_W223,MGM_W222);


	not MGM_G267(MGM_W225,SE$delay);


	and MGM_G268(ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE,MGM_W225,MGM_W224);


	not MGM_G269(MGM_W226,D2$delay);


	and MGM_G270(MGM_W227,MGM_W226,D1$delay);


	and MGM_G271(MGM_W228,SD$delay,MGM_W227);


	not MGM_G272(MGM_W229,SE$delay);


	and MGM_G273(ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE,MGM_W229,MGM_W228);


	not MGM_G274(MGM_W230,D1$delay);


	not MGM_G275(MGM_W231,D2$delay);


	and MGM_G276(MGM_W232,MGM_W231,MGM_W230);


	not MGM_G277(MGM_W233,S$delay);


	and MGM_G278(MGM_W234,MGM_W233,MGM_W232);


	and MGM_G279(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W234);


	not MGM_G280(MGM_W235,D1$delay);


	not MGM_G281(MGM_W236,D2$delay);


	and MGM_G282(MGM_W237,MGM_W236,MGM_W235);


	and MGM_G283(MGM_W238,S$delay,MGM_W237);


	and MGM_G284(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W238);


	not MGM_G285(MGM_W239,D1$delay);


	and MGM_G286(MGM_W240,D2$delay,MGM_W239);


	not MGM_G287(MGM_W241,S$delay);


	and MGM_G288(MGM_W242,MGM_W241,MGM_W240);


	and MGM_G289(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W242);


	not MGM_G290(MGM_W243,D1$delay);


	and MGM_G291(MGM_W244,D2$delay,MGM_W243);


	and MGM_G292(MGM_W245,S$delay,MGM_W244);


	and MGM_G293(ENABLE_NOT_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W245);


	not MGM_G294(MGM_W246,D2$delay);


	and MGM_G295(MGM_W247,MGM_W246,D1$delay);


	not MGM_G296(MGM_W248,S$delay);


	and MGM_G297(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G298(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W249);


	not MGM_G299(MGM_W250,D2$delay);


	and MGM_G300(MGM_W251,MGM_W250,D1$delay);


	and MGM_G301(MGM_W252,S$delay,MGM_W251);


	and MGM_G302(ENABLE_D1_AND_NOT_D2_AND_S_AND_SE,SE$delay,MGM_W252);


	and MGM_G303(MGM_W253,D2$delay,D1$delay);


	not MGM_G304(MGM_W254,S$delay);


	and MGM_G305(MGM_W255,MGM_W254,MGM_W253);


	and MGM_G306(ENABLE_D1_AND_D2_AND_NOT_S_AND_SE,SE$delay,MGM_W255);


	and MGM_G307(MGM_W256,D2$delay,D1$delay);


	and MGM_G308(MGM_W257,S$delay,MGM_W256);


	and MGM_G309(ENABLE_D1_AND_D2_AND_S_AND_SE,SE$delay,MGM_W257);


	not MGM_G310(MGM_W258,D1$delay);


	not MGM_G311(MGM_W259,D2$delay);


	and MGM_G312(MGM_W260,MGM_W259,MGM_W258);


	not MGM_G313(MGM_W261,S$delay);


	and MGM_G314(MGM_W262,MGM_W261,MGM_W260);


	and MGM_G315(ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W262);


	not MGM_G316(MGM_W263,D1$delay);


	not MGM_G317(MGM_W264,D2$delay);


	and MGM_G318(MGM_W265,MGM_W264,MGM_W263);


	and MGM_G319(MGM_W266,S$delay,MGM_W265);


	and MGM_G320(ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD,SD$delay,MGM_W266);


	not MGM_G321(MGM_W267,D1$delay);


	and MGM_G322(MGM_W268,D2$delay,MGM_W267);


	not MGM_G323(MGM_W269,S$delay);


	and MGM_G324(MGM_W270,MGM_W269,MGM_W268);


	not MGM_G325(MGM_W271,SD$delay);


	and MGM_G326(ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W271,MGM_W270);


	not MGM_G327(MGM_W272,D1$delay);


	and MGM_G328(MGM_W273,D2$delay,MGM_W272);


	and MGM_G329(MGM_W274,S$delay,MGM_W273);


	and MGM_G330(ENABLE_NOT_D1_AND_D2_AND_S_AND_SD,SD$delay,MGM_W274);


	not MGM_G331(MGM_W275,D2$delay);


	and MGM_G332(MGM_W276,MGM_W275,D1$delay);


	not MGM_G333(MGM_W277,S$delay);


	and MGM_G334(MGM_W278,MGM_W277,MGM_W276);


	and MGM_G335(ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD,SD$delay,MGM_W278);


	not MGM_G336(MGM_W279,D2$delay);


	and MGM_G337(MGM_W280,MGM_W279,D1$delay);


	and MGM_G338(MGM_W281,S$delay,MGM_W280);


	not MGM_G339(MGM_W282,SD$delay);


	and MGM_G340(ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD,MGM_W282,MGM_W281);


	and MGM_G341(MGM_W283,D2$delay,D1$delay);


	not MGM_G342(MGM_W284,S$delay);


	and MGM_G343(MGM_W285,MGM_W284,MGM_W283);


	not MGM_G344(MGM_W286,SD$delay);


	and MGM_G345(ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD,MGM_W286,MGM_W285);


	and MGM_G346(MGM_W287,D2$delay,D1$delay);


	and MGM_G347(MGM_W288,S$delay,MGM_W287);


	not MGM_G348(MGM_W289,SD$delay);


	and MGM_G349(ENABLE_D1_AND_D2_AND_S_AND_NOT_SD,MGM_W289,MGM_W288);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_NOT_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_D2_AND_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_D1_AND_NOT_S_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_D1_AND_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_D1_AND_NOT_D2_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D1_AND_D2_AND_S_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_NOT_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D1_AND_D2_AND_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_NOT_S_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_NOT_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_NOT_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D1_AND_D2_AND_S_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQM1HM( Q, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQM1HM_func SDFQM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQM1HM_func SDFQM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQM2HM( Q, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQM2HM_func SDFQM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQM2HM_func SDFQM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQM4HM( Q, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQM4HM_func SDFQM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQM4HM_func SDFQM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQM8HM( Q, CK, D, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQM8HM_func SDFQM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQM8HM_func SDFQM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,SD$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SE$delay);


	and MGM_G4(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W4,D$delay);


	not MGM_G6(MGM_W5,SD$delay);


	and MGM_G7(MGM_W6,MGM_W5,MGM_W4);


	and MGM_G8(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W6);


	not MGM_G9(MGM_W7,D$delay);


	and MGM_G10(MGM_W8,SD$delay,MGM_W7);


	not MGM_G11(MGM_W9,SE$delay);


	and MGM_G12(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W9,MGM_W8);


	not MGM_G13(MGM_W10,D$delay);


	and MGM_G14(MGM_W11,SD$delay,MGM_W10);


	and MGM_G15(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W11);


	not MGM_G16(MGM_W12,SD$delay);


	and MGM_G17(MGM_W13,MGM_W12,D$delay);


	not MGM_G18(MGM_W14,SE$delay);


	and MGM_G19(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W14,MGM_W13);


	not MGM_G20(MGM_W15,SD$delay);


	and MGM_G21(MGM_W16,MGM_W15,D$delay);


	and MGM_G22(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W16);


	and MGM_G23(MGM_W17,SD$delay,D$delay);


	not MGM_G24(MGM_W18,SE$delay);


	and MGM_G25(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W18,MGM_W17);


	and MGM_G26(MGM_W19,SD$delay,D$delay);


	and MGM_G27(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G28(MGM_W20,SD$delay);


	not MGM_G29(MGM_W21,SE$delay);


	and MGM_G30(ENABLE_NOT_SD_AND_NOT_SE,MGM_W21,MGM_W20);


	not MGM_G31(MGM_W22,SE$delay);


	and MGM_G32(ENABLE_SD_AND_NOT_SE,MGM_W22,SD$delay);


	not MGM_G33(MGM_W23,D$delay);


	and MGM_G34(ENABLE_NOT_D_AND_SE,SE$delay,MGM_W23);


	and MGM_G35(ENABLE_D_AND_SE,SE$delay,D$delay);


	not MGM_G36(MGM_W24,D$delay);


	and MGM_G37(ENABLE_NOT_D_AND_SD,SD$delay,MGM_W24);


	not MGM_G38(MGM_W25,SD$delay);


	and MGM_G39(ENABLE_D_AND_NOT_SD,MGM_W25,D$delay);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRM1HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRM1HM_func SDFQRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRM1HM_func SDFQRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRM2HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRM2HM_func SDFQRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRM2HM_func SDFQRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRM4HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRM4HM_func SDFQRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRM4HM_func SDFQRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRM8HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRM8HM_func SDFQRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRM8HM_func SDFQRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRSM1HM( Q, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM1HM_func SDFQRSM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRSM1HM_func SDFQRSM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRSM2HM( Q, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM2HM_func SDFQRSM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRSM2HM_func SDFQRSM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRSM4HM( Q, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM4HM_func SDFQRSM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRSM4HM_func SDFQRSM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRSM8HM( Q, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM8HM_func SDFQRSM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRSM8HM_func SDFQRSM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQRXM2HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQRXM2HM_func SDFQRXM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQRXM2HM_func SDFQRXM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQSM1HM( Q, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQSM1HM_func SDFQSM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQSM1HM_func SDFQSM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQSM2HM( Q, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQSM2HM_func SDFQSM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQSM2HM_func SDFQSM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQSM4HM( Q, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQSM4HM_func SDFQSM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQSM4HM_func SDFQSM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQSM8HM( Q, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQSM8HM_func SDFQSM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQSM8HM_func SDFQSM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQZRM1HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM1HM_func SDFQZRM1HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQZRM1HM_func SDFQZRM1HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQZRM2HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM2HM_func SDFQZRM2HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQZRM2HM_func SDFQZRM2HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQZRM4HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM4HM_func SDFQZRM4HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQZRM4HM_func SDFQZRM4HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFQZRM8HM( Q, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM8HM_func SDFQZRM8HM_behav_inst(.Q(Q),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFQZRM8HM_func SDFQZRM8HM_inst(.Q(Q),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRM1HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRM1HM_func SDFRM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRM1HM_func SDFRM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRM2HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRM2HM_func SDFRM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRM2HM_func SDFRM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRM4HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRM4HM_func SDFRM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRM4HM_func SDFRM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRM8HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRM8HM_func SDFRM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRM8HM_func SDFRM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,RB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,RB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,RB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,RB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,RB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,RB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,RB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,RB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,RB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	and MGM_G44(MGM_W34,SD$delay,MGM_W33);


	and MGM_G45(ENABLE_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W34);


	not MGM_G46(MGM_W35,SD$delay);


	and MGM_G47(MGM_W36,MGM_W35,D$delay);


	not MGM_G48(MGM_W37,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W37,MGM_W36);


	and MGM_G50(MGM_W38,SD$delay,D$delay);


	not MGM_G51(MGM_W39,SE$delay);


	and MGM_G52(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G53(MGM_W40,SD$delay,D$delay);


	and MGM_G54(ENABLE_D_AND_SD_AND_SE,SE$delay,MGM_W40);


	not MGM_G55(MGM_W41,CK$delay);


	not MGM_G56(MGM_W42,D$delay);


	and MGM_G57(MGM_W43,MGM_W42,MGM_W41);


	not MGM_G58(MGM_W44,SD$delay);


	and MGM_G59(MGM_W45,MGM_W44,MGM_W43);


	not MGM_G60(MGM_W46,SE$delay);


	and MGM_G61(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W47,CK$delay);


	not MGM_G63(MGM_W48,D$delay);


	and MGM_G64(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G65(MGM_W50,SD$delay);


	and MGM_G66(MGM_W51,MGM_W50,MGM_W49);


	and MGM_G67(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W51);


	not MGM_G68(MGM_W52,CK$delay);


	not MGM_G69(MGM_W53,D$delay);


	and MGM_G70(MGM_W54,MGM_W53,MGM_W52);


	and MGM_G71(MGM_W55,SD$delay,MGM_W54);


	not MGM_G72(MGM_W56,SE$delay);


	and MGM_G73(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W56,MGM_W55);


	not MGM_G74(MGM_W57,CK$delay);


	not MGM_G75(MGM_W58,D$delay);


	and MGM_G76(MGM_W59,MGM_W58,MGM_W57);


	and MGM_G77(MGM_W60,SD$delay,MGM_W59);


	and MGM_G78(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W60);


	not MGM_G79(MGM_W61,CK$delay);


	and MGM_G80(MGM_W62,D$delay,MGM_W61);


	not MGM_G81(MGM_W63,SD$delay);


	and MGM_G82(MGM_W64,MGM_W63,MGM_W62);


	not MGM_G83(MGM_W65,SE$delay);


	and MGM_G84(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W65,MGM_W64);


	not MGM_G85(MGM_W66,CK$delay);


	and MGM_G86(MGM_W67,D$delay,MGM_W66);


	not MGM_G87(MGM_W68,SD$delay);


	and MGM_G88(MGM_W69,MGM_W68,MGM_W67);


	and MGM_G89(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W69);


	not MGM_G90(MGM_W70,CK$delay);


	and MGM_G91(MGM_W71,D$delay,MGM_W70);


	and MGM_G92(MGM_W72,SD$delay,MGM_W71);


	not MGM_G93(MGM_W73,SE$delay);


	and MGM_G94(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G95(MGM_W74,CK$delay);


	and MGM_G96(MGM_W75,D$delay,MGM_W74);


	and MGM_G97(MGM_W76,SD$delay,MGM_W75);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W76);


	not MGM_G99(MGM_W77,D$delay);


	and MGM_G100(MGM_W78,MGM_W77,CK$delay);


	not MGM_G101(MGM_W79,SD$delay);


	and MGM_G102(MGM_W80,MGM_W79,MGM_W78);


	not MGM_G103(MGM_W81,SE$delay);


	and MGM_G104(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W81,MGM_W80);


	not MGM_G105(MGM_W82,D$delay);


	and MGM_G106(MGM_W83,MGM_W82,CK$delay);


	not MGM_G107(MGM_W84,SD$delay);


	and MGM_G108(MGM_W85,MGM_W84,MGM_W83);


	and MGM_G109(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W85);


	not MGM_G110(MGM_W86,D$delay);


	and MGM_G111(MGM_W87,MGM_W86,CK$delay);


	and MGM_G112(MGM_W88,SD$delay,MGM_W87);


	not MGM_G113(MGM_W89,SE$delay);


	and MGM_G114(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W89,MGM_W88);


	not MGM_G115(MGM_W90,D$delay);


	and MGM_G116(MGM_W91,MGM_W90,CK$delay);


	and MGM_G117(MGM_W92,SD$delay,MGM_W91);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W92);


	and MGM_G119(MGM_W93,D$delay,CK$delay);


	not MGM_G120(MGM_W94,SD$delay);


	and MGM_G121(MGM_W95,MGM_W94,MGM_W93);


	not MGM_G122(MGM_W96,SE$delay);


	and MGM_G123(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W96,MGM_W95);


	and MGM_G124(MGM_W97,D$delay,CK$delay);


	not MGM_G125(MGM_W98,SD$delay);


	and MGM_G126(MGM_W99,MGM_W98,MGM_W97);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W99);


	and MGM_G128(MGM_W100,D$delay,CK$delay);


	and MGM_G129(MGM_W101,SD$delay,MGM_W100);


	not MGM_G130(MGM_W102,SE$delay);


	and MGM_G131(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W102,MGM_W101);


	and MGM_G132(MGM_W103,D$delay,CK$delay);


	and MGM_G133(MGM_W104,SD$delay,MGM_W103);


	and MGM_G134(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W104);


	not MGM_G135(MGM_W105,D$delay);


	and MGM_G136(MGM_W106,RB$delay,MGM_W105);


	and MGM_G137(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W106);


	and MGM_G138(MGM_W107,RB$delay,D$delay);


	and MGM_G139(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W107);


	not MGM_G140(MGM_W108,D$delay);


	and MGM_G141(MGM_W109,RB$delay,MGM_W108);


	and MGM_G142(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W109);


	and MGM_G143(MGM_W110,RB$delay,D$delay);


	not MGM_G144(MGM_W111,SD$delay);


	and MGM_G145(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W111,MGM_W110);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRSM1HM( Q, QB, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRSM1HM_func SDFRSM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRSM1HM_func SDFRSM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRSM2HM( Q, QB, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRSM2HM_func SDFRSM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRSM2HM_func SDFRSM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRSM4HM( Q, QB, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRSM4HM_func SDFRSM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRSM4HM_func SDFRSM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFRSM8HM( Q, QB, CK, D, RB, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFRSM8HM_func SDFRSM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFRSM8HM_func SDFRSM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,RB$delay,MGM_W0);


	and MGM_G2(MGM_W2,SB$delay,MGM_W1);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	and MGM_G8(MGM_W7,RB$delay,MGM_W6);


	and MGM_G9(MGM_W8,SB$delay,MGM_W7);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	and MGM_G14(MGM_W12,RB$delay,MGM_W11);


	and MGM_G15(MGM_W13,SB$delay,MGM_W12);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	and MGM_G20(MGM_W17,RB$delay,MGM_W16);


	and MGM_G21(MGM_W18,SB$delay,MGM_W17);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W19);


	and MGM_G24(MGM_W20,RB$delay,D$delay);


	and MGM_G25(MGM_W21,SB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	and MGM_G30(MGM_W25,RB$delay,D$delay);


	and MGM_G31(MGM_W26,SB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	and MGM_G35(MGM_W29,RB$delay,D$delay);


	and MGM_G36(MGM_W30,SB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	and MGM_G40(MGM_W33,RB$delay,D$delay);


	and MGM_G41(MGM_W34,SB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W35);


	and MGM_G44(MGM_W36,SB$delay,RB$delay);


	not MGM_G45(MGM_W37,SD$delay);


	and MGM_G46(MGM_W38,MGM_W37,MGM_W36);


	not MGM_G47(MGM_W39,SE$delay);


	and MGM_G48(ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W39,MGM_W38);


	and MGM_G49(MGM_W40,SB$delay,RB$delay);


	and MGM_G50(MGM_W41,SD$delay,MGM_W40);


	not MGM_G51(MGM_W42,SE$delay);


	and MGM_G52(ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G53(MGM_W43,D$delay);


	and MGM_G54(MGM_W44,SB$delay,MGM_W43);


	and MGM_G55(MGM_W45,SD$delay,MGM_W44);


	and MGM_G56(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W45);


	and MGM_G57(MGM_W46,SB$delay,D$delay);


	not MGM_G58(MGM_W47,SD$delay);


	and MGM_G59(MGM_W48,MGM_W47,MGM_W46);


	not MGM_G60(MGM_W49,SE$delay);


	and MGM_G61(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W49,MGM_W48);


	and MGM_G62(MGM_W50,SB$delay,D$delay);


	and MGM_G63(MGM_W51,SD$delay,MGM_W50);


	not MGM_G64(MGM_W52,SE$delay);


	and MGM_G65(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W52,MGM_W51);


	and MGM_G66(MGM_W53,SB$delay,D$delay);


	and MGM_G67(MGM_W54,SD$delay,MGM_W53);


	and MGM_G68(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W54);


	not MGM_G69(MGM_W55,CK$delay);


	not MGM_G70(MGM_W56,D$delay);


	and MGM_G71(MGM_W57,MGM_W56,MGM_W55);


	and MGM_G72(MGM_W58,SB$delay,MGM_W57);


	not MGM_G73(MGM_W59,SD$delay);


	and MGM_G74(MGM_W60,MGM_W59,MGM_W58);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	not MGM_G77(MGM_W62,CK$delay);


	not MGM_G78(MGM_W63,D$delay);


	and MGM_G79(MGM_W64,MGM_W63,MGM_W62);


	and MGM_G80(MGM_W65,SB$delay,MGM_W64);


	not MGM_G81(MGM_W66,SD$delay);


	and MGM_G82(MGM_W67,MGM_W66,MGM_W65);


	and MGM_G83(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W67);


	not MGM_G84(MGM_W68,CK$delay);


	not MGM_G85(MGM_W69,D$delay);


	and MGM_G86(MGM_W70,MGM_W69,MGM_W68);


	and MGM_G87(MGM_W71,SB$delay,MGM_W70);


	and MGM_G88(MGM_W72,SD$delay,MGM_W71);


	not MGM_G89(MGM_W73,SE$delay);


	and MGM_G90(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G91(MGM_W74,CK$delay);


	not MGM_G92(MGM_W75,D$delay);


	and MGM_G93(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G94(MGM_W77,SB$delay,MGM_W76);


	and MGM_G95(MGM_W78,SD$delay,MGM_W77);


	and MGM_G96(ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W78);


	not MGM_G97(MGM_W79,CK$delay);


	and MGM_G98(MGM_W80,D$delay,MGM_W79);


	and MGM_G99(MGM_W81,SB$delay,MGM_W80);


	not MGM_G100(MGM_W82,SD$delay);


	and MGM_G101(MGM_W83,MGM_W82,MGM_W81);


	not MGM_G102(MGM_W84,SE$delay);


	and MGM_G103(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W84,MGM_W83);


	not MGM_G104(MGM_W85,CK$delay);


	and MGM_G105(MGM_W86,D$delay,MGM_W85);


	and MGM_G106(MGM_W87,SB$delay,MGM_W86);


	not MGM_G107(MGM_W88,SD$delay);


	and MGM_G108(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G109(ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G110(MGM_W90,CK$delay);


	and MGM_G111(MGM_W91,D$delay,MGM_W90);


	and MGM_G112(MGM_W92,SB$delay,MGM_W91);


	and MGM_G113(MGM_W93,SD$delay,MGM_W92);


	not MGM_G114(MGM_W94,SE$delay);


	and MGM_G115(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W94,MGM_W93);


	not MGM_G116(MGM_W95,CK$delay);


	and MGM_G117(MGM_W96,D$delay,MGM_W95);


	and MGM_G118(MGM_W97,SB$delay,MGM_W96);


	and MGM_G119(MGM_W98,SD$delay,MGM_W97);


	and MGM_G120(ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W98);


	not MGM_G121(MGM_W99,D$delay);


	and MGM_G122(MGM_W100,MGM_W99,CK$delay);


	and MGM_G123(MGM_W101,SB$delay,MGM_W100);


	not MGM_G124(MGM_W102,SD$delay);


	and MGM_G125(MGM_W103,MGM_W102,MGM_W101);


	not MGM_G126(MGM_W104,SE$delay);


	and MGM_G127(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W104,MGM_W103);


	not MGM_G128(MGM_W105,D$delay);


	and MGM_G129(MGM_W106,MGM_W105,CK$delay);


	and MGM_G130(MGM_W107,SB$delay,MGM_W106);


	not MGM_G131(MGM_W108,SD$delay);


	and MGM_G132(MGM_W109,MGM_W108,MGM_W107);


	and MGM_G133(ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W109);


	not MGM_G134(MGM_W110,D$delay);


	and MGM_G135(MGM_W111,MGM_W110,CK$delay);


	and MGM_G136(MGM_W112,SB$delay,MGM_W111);


	and MGM_G137(MGM_W113,SD$delay,MGM_W112);


	not MGM_G138(MGM_W114,SE$delay);


	and MGM_G139(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W114,MGM_W113);


	not MGM_G140(MGM_W115,D$delay);


	and MGM_G141(MGM_W116,MGM_W115,CK$delay);


	and MGM_G142(MGM_W117,SB$delay,MGM_W116);


	and MGM_G143(MGM_W118,SD$delay,MGM_W117);


	and MGM_G144(ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W118);


	and MGM_G145(MGM_W119,D$delay,CK$delay);


	and MGM_G146(MGM_W120,SB$delay,MGM_W119);


	not MGM_G147(MGM_W121,SD$delay);


	and MGM_G148(MGM_W122,MGM_W121,MGM_W120);


	not MGM_G149(MGM_W123,SE$delay);


	and MGM_G150(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W123,MGM_W122);


	and MGM_G151(MGM_W124,D$delay,CK$delay);


	and MGM_G152(MGM_W125,SB$delay,MGM_W124);


	not MGM_G153(MGM_W126,SD$delay);


	and MGM_G154(MGM_W127,MGM_W126,MGM_W125);


	and MGM_G155(ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W127);


	and MGM_G156(MGM_W128,D$delay,CK$delay);


	and MGM_G157(MGM_W129,SB$delay,MGM_W128);


	and MGM_G158(MGM_W130,SD$delay,MGM_W129);


	not MGM_G159(MGM_W131,SE$delay);


	and MGM_G160(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W131,MGM_W130);


	and MGM_G161(MGM_W132,D$delay,CK$delay);


	and MGM_G162(MGM_W133,SB$delay,MGM_W132);


	and MGM_G163(MGM_W134,SD$delay,MGM_W133);


	and MGM_G164(ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W134);


	not MGM_G165(MGM_W135,CK$delay);


	not MGM_G166(MGM_W136,D$delay);


	and MGM_G167(MGM_W137,MGM_W136,MGM_W135);


	not MGM_G168(MGM_W138,SD$delay);


	and MGM_G169(MGM_W139,MGM_W138,MGM_W137);


	not MGM_G170(MGM_W140,SE$delay);


	and MGM_G171(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W140,MGM_W139);


	not MGM_G172(MGM_W141,CK$delay);


	not MGM_G173(MGM_W142,D$delay);


	and MGM_G174(MGM_W143,MGM_W142,MGM_W141);


	not MGM_G175(MGM_W144,SD$delay);


	and MGM_G176(MGM_W145,MGM_W144,MGM_W143);


	and MGM_G177(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W145);


	not MGM_G178(MGM_W146,CK$delay);


	not MGM_G179(MGM_W147,D$delay);


	and MGM_G180(MGM_W148,MGM_W147,MGM_W146);


	and MGM_G181(MGM_W149,SD$delay,MGM_W148);


	not MGM_G182(MGM_W150,SE$delay);


	and MGM_G183(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W150,MGM_W149);


	not MGM_G184(MGM_W151,CK$delay);


	not MGM_G185(MGM_W152,D$delay);


	and MGM_G186(MGM_W153,MGM_W152,MGM_W151);


	and MGM_G187(MGM_W154,SD$delay,MGM_W153);


	and MGM_G188(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W154);


	not MGM_G189(MGM_W155,CK$delay);


	and MGM_G190(MGM_W156,D$delay,MGM_W155);


	not MGM_G191(MGM_W157,SD$delay);


	and MGM_G192(MGM_W158,MGM_W157,MGM_W156);


	not MGM_G193(MGM_W159,SE$delay);


	and MGM_G194(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W159,MGM_W158);


	not MGM_G195(MGM_W160,CK$delay);


	and MGM_G196(MGM_W161,D$delay,MGM_W160);


	not MGM_G197(MGM_W162,SD$delay);


	and MGM_G198(MGM_W163,MGM_W162,MGM_W161);


	and MGM_G199(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W163);


	not MGM_G200(MGM_W164,CK$delay);


	and MGM_G201(MGM_W165,D$delay,MGM_W164);


	and MGM_G202(MGM_W166,SD$delay,MGM_W165);


	not MGM_G203(MGM_W167,SE$delay);


	and MGM_G204(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W167,MGM_W166);


	not MGM_G205(MGM_W168,CK$delay);


	and MGM_G206(MGM_W169,D$delay,MGM_W168);


	and MGM_G207(MGM_W170,SD$delay,MGM_W169);


	and MGM_G208(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W170);


	not MGM_G209(MGM_W171,D$delay);


	and MGM_G210(MGM_W172,MGM_W171,CK$delay);


	not MGM_G211(MGM_W173,SD$delay);


	and MGM_G212(MGM_W174,MGM_W173,MGM_W172);


	not MGM_G213(MGM_W175,SE$delay);


	and MGM_G214(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W175,MGM_W174);


	not MGM_G215(MGM_W176,D$delay);


	and MGM_G216(MGM_W177,MGM_W176,CK$delay);


	not MGM_G217(MGM_W178,SD$delay);


	and MGM_G218(MGM_W179,MGM_W178,MGM_W177);


	and MGM_G219(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W179);


	not MGM_G220(MGM_W180,D$delay);


	and MGM_G221(MGM_W181,MGM_W180,CK$delay);


	and MGM_G222(MGM_W182,SD$delay,MGM_W181);


	not MGM_G223(MGM_W183,SE$delay);


	and MGM_G224(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W183,MGM_W182);


	not MGM_G225(MGM_W184,D$delay);


	and MGM_G226(MGM_W185,MGM_W184,CK$delay);


	and MGM_G227(MGM_W186,SD$delay,MGM_W185);


	and MGM_G228(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W186);


	and MGM_G229(MGM_W187,D$delay,CK$delay);


	not MGM_G230(MGM_W188,SD$delay);


	and MGM_G231(MGM_W189,MGM_W188,MGM_W187);


	not MGM_G232(MGM_W190,SE$delay);


	and MGM_G233(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W190,MGM_W189);


	and MGM_G234(MGM_W191,D$delay,CK$delay);


	not MGM_G235(MGM_W192,SD$delay);


	and MGM_G236(MGM_W193,MGM_W192,MGM_W191);


	and MGM_G237(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W193);


	and MGM_G238(MGM_W194,D$delay,CK$delay);


	and MGM_G239(MGM_W195,SD$delay,MGM_W194);


	not MGM_G240(MGM_W196,SE$delay);


	and MGM_G241(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W196,MGM_W195);


	and MGM_G242(MGM_W197,D$delay,CK$delay);


	and MGM_G243(MGM_W198,SD$delay,MGM_W197);


	and MGM_G244(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W198);


	not MGM_G245(MGM_W199,D$delay);


	and MGM_G246(MGM_W200,RB$delay,MGM_W199);


	not MGM_G247(MGM_W201,SD$delay);


	and MGM_G248(MGM_W202,MGM_W201,MGM_W200);


	not MGM_G249(MGM_W203,SE$delay);


	and MGM_G250(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W203,MGM_W202);


	not MGM_G251(MGM_W204,D$delay);


	and MGM_G252(MGM_W205,RB$delay,MGM_W204);


	not MGM_G253(MGM_W206,SD$delay);


	and MGM_G254(MGM_W207,MGM_W206,MGM_W205);


	and MGM_G255(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W207);


	not MGM_G256(MGM_W208,D$delay);


	and MGM_G257(MGM_W209,RB$delay,MGM_W208);


	and MGM_G258(MGM_W210,SD$delay,MGM_W209);


	not MGM_G259(MGM_W211,SE$delay);


	and MGM_G260(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W211,MGM_W210);


	and MGM_G261(MGM_W212,RB$delay,D$delay);


	not MGM_G262(MGM_W213,SD$delay);


	and MGM_G263(MGM_W214,MGM_W213,MGM_W212);


	and MGM_G264(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W214);


	not MGM_G265(MGM_W215,CK$delay);


	not MGM_G266(MGM_W216,D$delay);


	and MGM_G267(MGM_W217,MGM_W216,MGM_W215);


	and MGM_G268(MGM_W218,RB$delay,MGM_W217);


	not MGM_G269(MGM_W219,SD$delay);


	and MGM_G270(MGM_W220,MGM_W219,MGM_W218);


	not MGM_G271(MGM_W221,SE$delay);


	and MGM_G272(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W221,MGM_W220);


	not MGM_G273(MGM_W222,CK$delay);


	not MGM_G274(MGM_W223,D$delay);


	and MGM_G275(MGM_W224,MGM_W223,MGM_W222);


	and MGM_G276(MGM_W225,RB$delay,MGM_W224);


	not MGM_G277(MGM_W226,SD$delay);


	and MGM_G278(MGM_W227,MGM_W226,MGM_W225);


	and MGM_G279(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W227);


	not MGM_G280(MGM_W228,CK$delay);


	not MGM_G281(MGM_W229,D$delay);


	and MGM_G282(MGM_W230,MGM_W229,MGM_W228);


	and MGM_G283(MGM_W231,RB$delay,MGM_W230);


	and MGM_G284(MGM_W232,SD$delay,MGM_W231);


	not MGM_G285(MGM_W233,SE$delay);


	and MGM_G286(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W233,MGM_W232);


	not MGM_G287(MGM_W234,CK$delay);


	not MGM_G288(MGM_W235,D$delay);


	and MGM_G289(MGM_W236,MGM_W235,MGM_W234);


	and MGM_G290(MGM_W237,RB$delay,MGM_W236);


	and MGM_G291(MGM_W238,SD$delay,MGM_W237);


	and MGM_G292(ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W238);


	not MGM_G293(MGM_W239,CK$delay);


	and MGM_G294(MGM_W240,D$delay,MGM_W239);


	and MGM_G295(MGM_W241,RB$delay,MGM_W240);


	not MGM_G296(MGM_W242,SD$delay);


	and MGM_G297(MGM_W243,MGM_W242,MGM_W241);


	not MGM_G298(MGM_W244,SE$delay);


	and MGM_G299(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W244,MGM_W243);


	not MGM_G300(MGM_W245,CK$delay);


	and MGM_G301(MGM_W246,D$delay,MGM_W245);


	and MGM_G302(MGM_W247,RB$delay,MGM_W246);


	not MGM_G303(MGM_W248,SD$delay);


	and MGM_G304(MGM_W249,MGM_W248,MGM_W247);


	and MGM_G305(ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W249);


	not MGM_G306(MGM_W250,CK$delay);


	and MGM_G307(MGM_W251,D$delay,MGM_W250);


	and MGM_G308(MGM_W252,RB$delay,MGM_W251);


	and MGM_G309(MGM_W253,SD$delay,MGM_W252);


	not MGM_G310(MGM_W254,SE$delay);


	and MGM_G311(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W254,MGM_W253);


	not MGM_G312(MGM_W255,CK$delay);


	and MGM_G313(MGM_W256,D$delay,MGM_W255);


	and MGM_G314(MGM_W257,RB$delay,MGM_W256);


	and MGM_G315(MGM_W258,SD$delay,MGM_W257);


	and MGM_G316(ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W258);


	not MGM_G317(MGM_W259,D$delay);


	and MGM_G318(MGM_W260,MGM_W259,CK$delay);


	and MGM_G319(MGM_W261,RB$delay,MGM_W260);


	not MGM_G320(MGM_W262,SD$delay);


	and MGM_G321(MGM_W263,MGM_W262,MGM_W261);


	not MGM_G322(MGM_W264,SE$delay);


	and MGM_G323(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W264,MGM_W263);


	not MGM_G324(MGM_W265,D$delay);


	and MGM_G325(MGM_W266,MGM_W265,CK$delay);


	and MGM_G326(MGM_W267,RB$delay,MGM_W266);


	not MGM_G327(MGM_W268,SD$delay);


	and MGM_G328(MGM_W269,MGM_W268,MGM_W267);


	and MGM_G329(ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W269);


	not MGM_G330(MGM_W270,D$delay);


	and MGM_G331(MGM_W271,MGM_W270,CK$delay);


	and MGM_G332(MGM_W272,RB$delay,MGM_W271);


	and MGM_G333(MGM_W273,SD$delay,MGM_W272);


	not MGM_G334(MGM_W274,SE$delay);


	and MGM_G335(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W274,MGM_W273);


	not MGM_G336(MGM_W275,D$delay);


	and MGM_G337(MGM_W276,MGM_W275,CK$delay);


	and MGM_G338(MGM_W277,RB$delay,MGM_W276);


	and MGM_G339(MGM_W278,SD$delay,MGM_W277);


	and MGM_G340(ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W278);


	and MGM_G341(MGM_W279,D$delay,CK$delay);


	and MGM_G342(MGM_W280,RB$delay,MGM_W279);


	not MGM_G343(MGM_W281,SD$delay);


	and MGM_G344(MGM_W282,MGM_W281,MGM_W280);


	not MGM_G345(MGM_W283,SE$delay);


	and MGM_G346(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W283,MGM_W282);


	and MGM_G347(MGM_W284,D$delay,CK$delay);


	and MGM_G348(MGM_W285,RB$delay,MGM_W284);


	not MGM_G349(MGM_W286,SD$delay);


	and MGM_G350(MGM_W287,MGM_W286,MGM_W285);


	and MGM_G351(ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W287);


	and MGM_G352(MGM_W288,D$delay,CK$delay);


	and MGM_G353(MGM_W289,RB$delay,MGM_W288);


	and MGM_G354(MGM_W290,SD$delay,MGM_W289);


	not MGM_G355(MGM_W291,SE$delay);


	and MGM_G356(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W291,MGM_W290);


	and MGM_G357(MGM_W292,D$delay,CK$delay);


	and MGM_G358(MGM_W293,RB$delay,MGM_W292);


	and MGM_G359(MGM_W294,SD$delay,MGM_W293);


	and MGM_G360(ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W294);


	not MGM_G361(MGM_W295,D$delay);


	and MGM_G362(MGM_W296,RB$delay,MGM_W295);


	and MGM_G363(MGM_W297,SB$delay,MGM_W296);


	and MGM_G364(ENABLE_NOT_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W297);


	and MGM_G365(MGM_W298,RB$delay,D$delay);


	and MGM_G366(MGM_W299,SB$delay,MGM_W298);


	and MGM_G367(ENABLE_D_AND_RB_AND_SB_AND_SE,SE$delay,MGM_W299);


	not MGM_G368(MGM_W300,D$delay);


	and MGM_G369(MGM_W301,RB$delay,MGM_W300);


	and MGM_G370(MGM_W302,SB$delay,MGM_W301);


	and MGM_G371(ENABLE_NOT_D_AND_RB_AND_SB_AND_SD,SD$delay,MGM_W302);


	and MGM_G372(MGM_W303,RB$delay,D$delay);


	and MGM_G373(MGM_W304,SB$delay,MGM_W303);


	not MGM_G374(MGM_W305,SD$delay);


	and MGM_G375(ENABLE_D_AND_RB_AND_SB_AND_NOT_SD,MGM_W305,MGM_W304);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge RB &&& (ENABLE_CK_AND_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// setuphold RB- SB-LH
	$setuphold(posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,RB$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	// setuphold SB- RB-LH
	$setuphold(posedge RB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		posedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,RB$delay,SB$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw RB_hl 
	$width(negedge RB,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFSM1HM( Q, QB, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFSM1HM_func SDFSM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFSM1HM_func SDFSM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFSM2HM( Q, QB, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFSM2HM_func SDFSM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFSM2HM_func SDFSM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFSM4HM( Q, QB, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFSM4HM_func SDFSM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFSM4HM_func SDFSM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFSM8HM( Q, QB, CK, D, SB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFSM8HM_func SDFSM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire SB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFSM8HM_func SDFSM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	and MGM_G1(MGM_W1,SB$delay,MGM_W0);


	not MGM_G2(MGM_W2,SD$delay);


	and MGM_G3(MGM_W3,MGM_W2,MGM_W1);


	not MGM_G4(MGM_W4,SE$delay);


	and MGM_G5(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W4,MGM_W3);


	not MGM_G6(MGM_W5,D$delay);


	and MGM_G7(MGM_W6,SB$delay,MGM_W5);


	not MGM_G8(MGM_W7,SD$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	and MGM_G10(ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W8);


	not MGM_G11(MGM_W9,D$delay);


	and MGM_G12(MGM_W10,SB$delay,MGM_W9);


	and MGM_G13(MGM_W11,SD$delay,MGM_W10);


	not MGM_G14(MGM_W12,SE$delay);


	and MGM_G15(ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W12,MGM_W11);


	not MGM_G16(MGM_W13,D$delay);


	and MGM_G17(MGM_W14,SB$delay,MGM_W13);


	and MGM_G18(MGM_W15,SD$delay,MGM_W14);


	and MGM_G19(ENABLE_NOT_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W15);


	and MGM_G20(MGM_W16,SB$delay,D$delay);


	not MGM_G21(MGM_W17,SD$delay);


	and MGM_G22(MGM_W18,MGM_W17,MGM_W16);


	not MGM_G23(MGM_W19,SE$delay);


	and MGM_G24(ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE,MGM_W19,MGM_W18);


	and MGM_G25(MGM_W20,SB$delay,D$delay);


	not MGM_G26(MGM_W21,SD$delay);


	and MGM_G27(MGM_W22,MGM_W21,MGM_W20);


	and MGM_G28(ENABLE_D_AND_SB_AND_NOT_SD_AND_SE,SE$delay,MGM_W22);


	and MGM_G29(MGM_W23,SB$delay,D$delay);


	and MGM_G30(MGM_W24,SD$delay,MGM_W23);


	not MGM_G31(MGM_W25,SE$delay);


	and MGM_G32(ENABLE_D_AND_SB_AND_SD_AND_NOT_SE,MGM_W25,MGM_W24);


	and MGM_G33(MGM_W26,SB$delay,D$delay);


	and MGM_G34(MGM_W27,SD$delay,MGM_W26);


	and MGM_G35(ENABLE_D_AND_SB_AND_SD_AND_SE,SE$delay,MGM_W27);


	not MGM_G36(MGM_W28,SD$delay);


	and MGM_G37(MGM_W29,MGM_W28,SB$delay);


	not MGM_G38(MGM_W30,SE$delay);


	and MGM_G39(ENABLE_SB_AND_NOT_SD_AND_NOT_SE,MGM_W30,MGM_W29);


	and MGM_G40(MGM_W31,SD$delay,SB$delay);


	not MGM_G41(MGM_W32,SE$delay);


	and MGM_G42(ENABLE_SB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G43(MGM_W33,D$delay);


	not MGM_G44(MGM_W34,SD$delay);


	and MGM_G45(MGM_W35,MGM_W34,MGM_W33);


	not MGM_G46(MGM_W36,SE$delay);


	and MGM_G47(ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W36,MGM_W35);


	not MGM_G48(MGM_W37,D$delay);


	not MGM_G49(MGM_W38,SD$delay);


	and MGM_G50(MGM_W39,MGM_W38,MGM_W37);


	and MGM_G51(ENABLE_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W39);


	not MGM_G52(MGM_W40,D$delay);


	and MGM_G53(MGM_W41,SD$delay,MGM_W40);


	not MGM_G54(MGM_W42,SE$delay);


	and MGM_G55(ENABLE_NOT_D_AND_SD_AND_NOT_SE,MGM_W42,MGM_W41);


	not MGM_G56(MGM_W43,SD$delay);


	and MGM_G57(MGM_W44,MGM_W43,D$delay);


	and MGM_G58(ENABLE_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G59(MGM_W45,CK$delay);


	not MGM_G60(MGM_W46,D$delay);


	and MGM_G61(MGM_W47,MGM_W46,MGM_W45);


	not MGM_G62(MGM_W48,SD$delay);


	and MGM_G63(MGM_W49,MGM_W48,MGM_W47);


	not MGM_G64(MGM_W50,SE$delay);


	and MGM_G65(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W50,MGM_W49);


	not MGM_G66(MGM_W51,CK$delay);


	not MGM_G67(MGM_W52,D$delay);


	and MGM_G68(MGM_W53,MGM_W52,MGM_W51);


	not MGM_G69(MGM_W54,SD$delay);


	and MGM_G70(MGM_W55,MGM_W54,MGM_W53);


	and MGM_G71(ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W55);


	not MGM_G72(MGM_W56,CK$delay);


	not MGM_G73(MGM_W57,D$delay);


	and MGM_G74(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G75(MGM_W59,SD$delay,MGM_W58);


	not MGM_G76(MGM_W60,SE$delay);


	and MGM_G77(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W60,MGM_W59);


	not MGM_G78(MGM_W61,CK$delay);


	not MGM_G79(MGM_W62,D$delay);


	and MGM_G80(MGM_W63,MGM_W62,MGM_W61);


	and MGM_G81(MGM_W64,SD$delay,MGM_W63);


	and MGM_G82(ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W64);


	not MGM_G83(MGM_W65,CK$delay);


	and MGM_G84(MGM_W66,D$delay,MGM_W65);


	not MGM_G85(MGM_W67,SD$delay);


	and MGM_G86(MGM_W68,MGM_W67,MGM_W66);


	not MGM_G87(MGM_W69,SE$delay);


	and MGM_G88(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W69,MGM_W68);


	not MGM_G89(MGM_W70,CK$delay);


	and MGM_G90(MGM_W71,D$delay,MGM_W70);


	not MGM_G91(MGM_W72,SD$delay);


	and MGM_G92(MGM_W73,MGM_W72,MGM_W71);


	and MGM_G93(ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W73);


	not MGM_G94(MGM_W74,CK$delay);


	and MGM_G95(MGM_W75,D$delay,MGM_W74);


	and MGM_G96(MGM_W76,SD$delay,MGM_W75);


	not MGM_G97(MGM_W77,SE$delay);


	and MGM_G98(ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W77,MGM_W76);


	not MGM_G99(MGM_W78,CK$delay);


	and MGM_G100(MGM_W79,D$delay,MGM_W78);


	and MGM_G101(MGM_W80,SD$delay,MGM_W79);


	and MGM_G102(ENABLE_NOT_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W80);


	not MGM_G103(MGM_W81,D$delay);


	and MGM_G104(MGM_W82,MGM_W81,CK$delay);


	not MGM_G105(MGM_W83,SD$delay);


	and MGM_G106(MGM_W84,MGM_W83,MGM_W82);


	not MGM_G107(MGM_W85,SE$delay);


	and MGM_G108(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE,MGM_W85,MGM_W84);


	not MGM_G109(MGM_W86,D$delay);


	and MGM_G110(MGM_W87,MGM_W86,CK$delay);


	not MGM_G111(MGM_W88,SD$delay);


	and MGM_G112(MGM_W89,MGM_W88,MGM_W87);


	and MGM_G113(ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W89);


	not MGM_G114(MGM_W90,D$delay);


	and MGM_G115(MGM_W91,MGM_W90,CK$delay);


	and MGM_G116(MGM_W92,SD$delay,MGM_W91);


	not MGM_G117(MGM_W93,SE$delay);


	and MGM_G118(ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE,MGM_W93,MGM_W92);


	not MGM_G119(MGM_W94,D$delay);


	and MGM_G120(MGM_W95,MGM_W94,CK$delay);


	and MGM_G121(MGM_W96,SD$delay,MGM_W95);


	and MGM_G122(ENABLE_CK_AND_NOT_D_AND_SD_AND_SE,SE$delay,MGM_W96);


	and MGM_G123(MGM_W97,D$delay,CK$delay);


	not MGM_G124(MGM_W98,SD$delay);


	and MGM_G125(MGM_W99,MGM_W98,MGM_W97);


	not MGM_G126(MGM_W100,SE$delay);


	and MGM_G127(ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE,MGM_W100,MGM_W99);


	and MGM_G128(MGM_W101,D$delay,CK$delay);


	not MGM_G129(MGM_W102,SD$delay);


	and MGM_G130(MGM_W103,MGM_W102,MGM_W101);


	and MGM_G131(ENABLE_CK_AND_D_AND_NOT_SD_AND_SE,SE$delay,MGM_W103);


	and MGM_G132(MGM_W104,D$delay,CK$delay);


	and MGM_G133(MGM_W105,SD$delay,MGM_W104);


	not MGM_G134(MGM_W106,SE$delay);


	and MGM_G135(ENABLE_CK_AND_D_AND_SD_AND_NOT_SE,MGM_W106,MGM_W105);


	and MGM_G136(MGM_W107,D$delay,CK$delay);


	and MGM_G137(MGM_W108,SD$delay,MGM_W107);


	and MGM_G138(ENABLE_CK_AND_D_AND_SD_AND_SE,SE$delay,MGM_W108);


	not MGM_G139(MGM_W109,D$delay);


	and MGM_G140(MGM_W110,SB$delay,MGM_W109);


	and MGM_G141(ENABLE_NOT_D_AND_SB_AND_SE,SE$delay,MGM_W110);


	and MGM_G142(MGM_W111,SB$delay,D$delay);


	and MGM_G143(ENABLE_D_AND_SB_AND_SE,SE$delay,MGM_W111);


	not MGM_G144(MGM_W112,D$delay);


	and MGM_G145(MGM_W113,SB$delay,MGM_W112);


	and MGM_G146(ENABLE_NOT_D_AND_SB_AND_SD,SD$delay,MGM_W113);


	and MGM_G147(MGM_W114,SB$delay,D$delay);


	not MGM_G148(MGM_W115,SD$delay);


	and MGM_G149(ENABLE_D_AND_SB_AND_NOT_SD,MGM_W115,MGM_W114);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// seq arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_SB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge CK &&& (ENABLE_NOT_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_SE === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_NOT_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_NOT_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge SB &&& (ENABLE_CK_AND_D_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_SB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_SB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// mpw SB_hl 
	$width(negedge SB,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFZRM1HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFZRM1HM_func SDFZRM1HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFZRM1HM_func SDFZRM1HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFZRM2HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFZRM2HM_func SDFZRM2HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFZRM2HM_func SDFZRM2HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFZRM4HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFZRM4HM_func SDFZRM4HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFZRM4HM_func SDFZRM4HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module SDFZRM8HM( Q, QB, CK, D, RB, SD, SE , VDD, VSS);
inout VDD;
inout VSS;
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

	SDFZRM8HM_func SDFZRM8HM_behav_inst(.Q(Q),.QB(QB),.CK(CK),.D(D),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier),.VDD(VDD),.VSS(VSS));

   `else

	wire CK$delay ;

	wire D$delay ;

	wire RB$delay ;

	wire SD$delay ;

	wire SE$delay ;

	SDFZRM8HM_func SDFZRM8HM_inst(.Q(Q),.QB(QB),.CK(CK$delay),.D(D$delay),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	not MGM_G0(MGM_W0,D$delay);


	not MGM_G1(MGM_W1,RB$delay);


	and MGM_G2(MGM_W2,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W3,SD$delay);


	and MGM_G4(MGM_W4,MGM_W3,MGM_W2);


	not MGM_G5(MGM_W5,SE$delay);


	and MGM_G6(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W5,MGM_W4);


	not MGM_G7(MGM_W6,D$delay);


	not MGM_G8(MGM_W7,RB$delay);


	and MGM_G9(MGM_W8,MGM_W7,MGM_W6);


	not MGM_G10(MGM_W9,SD$delay);


	and MGM_G11(MGM_W10,MGM_W9,MGM_W8);


	and MGM_G12(ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W10);


	not MGM_G13(MGM_W11,D$delay);


	not MGM_G14(MGM_W12,RB$delay);


	and MGM_G15(MGM_W13,MGM_W12,MGM_W11);


	and MGM_G16(MGM_W14,SD$delay,MGM_W13);


	not MGM_G17(MGM_W15,SE$delay);


	and MGM_G18(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W15,MGM_W14);


	not MGM_G19(MGM_W16,D$delay);


	not MGM_G20(MGM_W17,RB$delay);


	and MGM_G21(MGM_W18,MGM_W17,MGM_W16);


	and MGM_G22(MGM_W19,SD$delay,MGM_W18);


	and MGM_G23(ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W19);


	not MGM_G24(MGM_W20,D$delay);


	and MGM_G25(MGM_W21,RB$delay,MGM_W20);


	not MGM_G26(MGM_W22,SD$delay);


	and MGM_G27(MGM_W23,MGM_W22,MGM_W21);


	not MGM_G28(MGM_W24,SE$delay);


	and MGM_G29(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W24,MGM_W23);


	not MGM_G30(MGM_W25,D$delay);


	and MGM_G31(MGM_W26,RB$delay,MGM_W25);


	not MGM_G32(MGM_W27,SD$delay);


	and MGM_G33(MGM_W28,MGM_W27,MGM_W26);


	and MGM_G34(ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W28);


	not MGM_G35(MGM_W29,D$delay);


	and MGM_G36(MGM_W30,RB$delay,MGM_W29);


	and MGM_G37(MGM_W31,SD$delay,MGM_W30);


	not MGM_G38(MGM_W32,SE$delay);


	and MGM_G39(ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W32,MGM_W31);


	not MGM_G40(MGM_W33,D$delay);


	and MGM_G41(MGM_W34,RB$delay,MGM_W33);


	and MGM_G42(MGM_W35,SD$delay,MGM_W34);


	and MGM_G43(ENABLE_NOT_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W35);


	not MGM_G44(MGM_W36,RB$delay);


	and MGM_G45(MGM_W37,MGM_W36,D$delay);


	not MGM_G46(MGM_W38,SD$delay);


	and MGM_G47(MGM_W39,MGM_W38,MGM_W37);


	not MGM_G48(MGM_W40,SE$delay);


	and MGM_G49(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE,MGM_W40,MGM_W39);


	not MGM_G50(MGM_W41,RB$delay);


	and MGM_G51(MGM_W42,MGM_W41,D$delay);


	not MGM_G52(MGM_W43,SD$delay);


	and MGM_G53(MGM_W44,MGM_W43,MGM_W42);


	and MGM_G54(ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W44);


	not MGM_G55(MGM_W45,RB$delay);


	and MGM_G56(MGM_W46,MGM_W45,D$delay);


	and MGM_G57(MGM_W47,SD$delay,MGM_W46);


	not MGM_G58(MGM_W48,SE$delay);


	and MGM_G59(ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE,MGM_W48,MGM_W47);


	not MGM_G60(MGM_W49,RB$delay);


	and MGM_G61(MGM_W50,MGM_W49,D$delay);


	and MGM_G62(MGM_W51,SD$delay,MGM_W50);


	and MGM_G63(ENABLE_D_AND_NOT_RB_AND_SD_AND_SE,SE$delay,MGM_W51);


	and MGM_G64(MGM_W52,RB$delay,D$delay);


	not MGM_G65(MGM_W53,SD$delay);


	and MGM_G66(MGM_W54,MGM_W53,MGM_W52);


	not MGM_G67(MGM_W55,SE$delay);


	and MGM_G68(ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE,MGM_W55,MGM_W54);


	and MGM_G69(MGM_W56,RB$delay,D$delay);


	not MGM_G70(MGM_W57,SD$delay);


	and MGM_G71(MGM_W58,MGM_W57,MGM_W56);


	and MGM_G72(ENABLE_D_AND_RB_AND_NOT_SD_AND_SE,SE$delay,MGM_W58);


	and MGM_G73(MGM_W59,RB$delay,D$delay);


	and MGM_G74(MGM_W60,SD$delay,MGM_W59);


	not MGM_G75(MGM_W61,SE$delay);


	and MGM_G76(ENABLE_D_AND_RB_AND_SD_AND_NOT_SE,MGM_W61,MGM_W60);


	and MGM_G77(MGM_W62,RB$delay,D$delay);


	and MGM_G78(MGM_W63,SD$delay,MGM_W62);


	and MGM_G79(ENABLE_D_AND_RB_AND_SD_AND_SE,SE$delay,MGM_W63);


	not MGM_G80(MGM_W64,SD$delay);


	and MGM_G81(MGM_W65,MGM_W64,RB$delay);


	not MGM_G82(MGM_W66,SE$delay);


	and MGM_G83(ENABLE_RB_AND_NOT_SD_AND_NOT_SE,MGM_W66,MGM_W65);


	and MGM_G84(MGM_W67,SD$delay,RB$delay);


	not MGM_G85(MGM_W68,SE$delay);


	and MGM_G86(ENABLE_RB_AND_SD_AND_NOT_SE,MGM_W68,MGM_W67);


	not MGM_G87(MGM_W69,SD$delay);


	and MGM_G88(MGM_W70,MGM_W69,D$delay);


	not MGM_G89(MGM_W71,SE$delay);


	and MGM_G90(ENABLE_D_AND_NOT_SD_AND_NOT_SE,MGM_W71,MGM_W70);


	and MGM_G91(MGM_W72,SD$delay,D$delay);


	not MGM_G92(MGM_W73,SE$delay);


	and MGM_G93(ENABLE_D_AND_SD_AND_NOT_SE,MGM_W73,MGM_W72);


	not MGM_G94(MGM_W74,D$delay);


	not MGM_G95(MGM_W75,RB$delay);


	and MGM_G96(MGM_W76,MGM_W75,MGM_W74);


	and MGM_G97(ENABLE_NOT_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W76);


	not MGM_G98(MGM_W77,D$delay);


	and MGM_G99(MGM_W78,RB$delay,MGM_W77);


	and MGM_G100(ENABLE_NOT_D_AND_RB_AND_SE,SE$delay,MGM_W78);


	not MGM_G101(MGM_W79,RB$delay);


	and MGM_G102(MGM_W80,MGM_W79,D$delay);


	and MGM_G103(ENABLE_D_AND_NOT_RB_AND_SE,SE$delay,MGM_W80);


	and MGM_G104(MGM_W81,RB$delay,D$delay);


	and MGM_G105(ENABLE_D_AND_RB_AND_SE,SE$delay,MGM_W81);


	not MGM_G106(MGM_W82,D$delay);


	not MGM_G107(MGM_W83,RB$delay);


	and MGM_G108(MGM_W84,MGM_W83,MGM_W82);


	and MGM_G109(ENABLE_NOT_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W84);


	not MGM_G110(MGM_W85,D$delay);


	and MGM_G111(MGM_W86,RB$delay,MGM_W85);


	and MGM_G112(ENABLE_NOT_D_AND_RB_AND_SD,SD$delay,MGM_W86);


	not MGM_G113(MGM_W87,RB$delay);


	and MGM_G114(MGM_W88,MGM_W87,D$delay);


	and MGM_G115(ENABLE_D_AND_NOT_RB_AND_SD,SD$delay,MGM_W88);


	and MGM_G116(MGM_W89,RB$delay,D$delay);


	not MGM_G117(MGM_W90,SD$delay);


	and MGM_G118(ENABLE_D_AND_RB_AND_NOT_SD,MGM_W90,MGM_W89);


	// spec_gates_end



   specify

	// specify_block_begin 

	// seq arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// seq arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_NOT_SE === 1'b1)
		,1.0,0,notifier);

	$width(negedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	$width(posedge CK &&& (ENABLE_D_AND_RB_AND_SD_AND_SE === 1'b1)
		,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_NOT_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_D_AND_SD_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_NOT_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_NOT_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_D_AND_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_NOT_D_AND_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_NOT_RB_AND_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		posedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		negedge SE &&& (ENABLE_D_AND_RB_AND_NOT_SD === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// mpw CK_lh 
	$width(posedge CK,1.0,0,notifier);

	// mpw CK_hl 
	$width(negedge CK,1.0,0,notifier);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module TIE0HM( Z , VDD, VSS);
inout VDD;
inout VSS;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	TIE0HM_func TIE0HM_behav_inst(.Z(Z),.VDD(VDD),.VSS(VSS));

   `else

	TIE0HM_func TIE0HM_inst(.Z(Z),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module TIE1HM( Z , VDD, VSS);
inout VDD;
inout VSS;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	TIE1HM_func TIE1HM_behav_inst(.Z(Z),.VDD(VDD),.VSS(VSS));

   `else

	TIE1HM_func TIE1HM_inst(.Z(Z),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR2M0HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR2M0HM_func XNR2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XNR2M0HM_func XNR2M0HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR2M1HM_func XNR2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XNR2M1HM_func XNR2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR2M2HM_func XNR2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XNR2M2HM_func XNR2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR2M4HM_func XNR2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XNR2M4HM_func XNR2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR3M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR3M0HM_func XNR3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XNR3M0HM_func XNR3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR3M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR3M1HM_func XNR3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XNR3M1HM_func XNR3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR3M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR3M2HM_func XNR3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XNR3M2HM_func XNR3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR3M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR3M4HM_func XNR3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XNR3M4HM_func XNR3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR4M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR4M0HM_func XNR4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XNR4M0HM_func XNR4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR4M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR4M1HM_func XNR4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XNR4M1HM_func XNR4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR4M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR4M2HM_func XNR4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XNR4M2HM_func XNR4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XNR4M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XNR4M4HM_func XNR4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XNR4M4HM_func XNR4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M0HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M0HM_func XOR2M0HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M0HM_func XOR2M0HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M1HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M1HM_func XOR2M1HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M1HM_func XOR2M1HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M2HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M2HM_func XOR2M2HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M2HM_func XOR2M2HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M3HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M3HM_func XOR2M3HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M3HM_func XOR2M3HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M4HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M4HM_func XOR2M4HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M4HM_func XOR2M4HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M6HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M6HM_func XOR2M6HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M6HM_func XOR2M6HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR2M8HM( Z, A, B , VDD, VSS);
inout VDD;
inout VSS;
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR2M8HM_func XOR2M8HM_behav_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));

   `else

	XOR2M8HM_func XOR2M8HM_inst(.Z(Z),.A(A),.B(B),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR3M0HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR3M0HM_func XOR3M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XOR3M0HM_func XOR3M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR3M1HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR3M1HM_func XOR3M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XOR3M1HM_func XOR3M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR3M2HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR3M2HM_func XOR3M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XOR3M2HM_func XOR3M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR3M4HM( Z, A, B, C , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR3M4HM_func XOR3M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));

   `else

	XOR3M4HM_func XOR3M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR4M0HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR4M0HM_func XOR4M0HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XOR4M0HM_func XOR4M0HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR4M1HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR4M1HM_func XOR4M1HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XOR4M1HM_func XOR4M1HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR4M2HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR4M2HM_func XOR4M2HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XOR4M2HM_func XOR4M2HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module XOR4M4HM( Z, A, B, C, D , VDD, VSS);
inout VDD;
inout VSS;
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

	XOR4M4HM_func XOR4M4HM_behav_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));

   `else

	XOR4M4HM_func XOR4M4HM_inst(.Z(Z),.A(A),.B(B),.C(C),.D(D),.VDD(VDD),.VSS(VSS));


	// spec_gates_begin


	// spec_gates_end



   specify

	// specify_block_begin 

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	ifnone
	// comb arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// comb arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	ifnone
	// comb arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// comb arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

	ifnone
	// comb arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// comb arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// comb arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

	ifnone
	// comb arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// comb arc D --> Z
	 (D => Z) = (1.0,1.0);

	// specify_block_end 

   endspecify

   `endif 

endmodule
`endcelldefine

`celldefine
module ADFM0HM_func( CO, S, A, B, CI, VDD , VSS );
inout VSS;
inout VDD;
input A, B, CI;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (CI_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CI_org, CI, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(CO,A_org,B_org,CI_org); 

	ADFCSIOM2HM_udp_0(S,A_org,B_org,CI_org); 
endmodule
`endcelldefine

`celldefine
module ADFM1HM_func( CO, S, A, B, CI, VDD , VSS );
inout VSS;
inout VDD;
input A, B, CI;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (CI_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CI_org, CI, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(CO,A_org,B_org,CI_org); 

	ADFCSIOM2HM_udp_0(S,A_org,B_org,CI_org); 
endmodule
`endcelldefine

`celldefine
module ADFM2HM_func( CO, S, A, B, CI, VDD , VSS );
inout VSS;
inout VDD;
input A, B, CI;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (CI_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CI_org, CI, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(CO,A_org,B_org,CI_org); 

	ADFCSIOM2HM_udp_0(S,A_org,B_org,CI_org); 
endmodule
`endcelldefine

`celldefine
module ADFM4HM_func( CO, S, A, B, CI, VDD , VSS );
inout VSS;
inout VDD;
input A, B, CI;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (CI_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CI_org, CI, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(CO,A_org,B_org,CI_org); 

	ADFCSIOM2HM_udp_0(S,A_org,B_org,CI_org); 
endmodule
`endcelldefine

`celldefine
module ADFM8HM_func( CO, S, A, B, CI, VDD , VSS );
inout VSS;
inout VDD;
input A, B, CI;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (CI_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CI_org, CI, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(CO,A_org,B_org,CI_org); 

	ADFCSIOM2HM_udp_0(S,A_org,B_org,CI_org); 
endmodule
`endcelldefine

`celldefine
module ADHM0HM_func( CO, S, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(CO,A_org,B_org); 

	ADHM1HM_udp_1(S,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ADHM1HM_func( CO, S, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(CO,A_org,B_org); 

	ADHM1HM_udp_1(S,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ADHM2HM_func( CO, S, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(CO,A_org,B_org); 

	ADHM1HM_udp_1(S,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ADHM4HM_func( CO, S, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(CO,A_org,B_org); 

	ADHM1HM_udp_1(S,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ADHM8HM_func( CO, S, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output CO, S;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(CO,A_org,B_org); 

	ADHM1HM_udp_1(S,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M0HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M16HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AN3M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M12HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M16HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M6HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN3M8HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AN4M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M12HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M16HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M6HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AN4M8HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AN4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module AO211M0HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO211M1HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO211M1HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO211M1HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO211M2HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO211M1HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO211M4HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO211M1HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO211M8HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO211M1HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO21M0HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO21M1HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO21M2HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO21M4HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO21M8HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO221M0HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO221M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO221M1HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO221M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO221M2HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO221M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO221M4HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO221M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO221M8HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO221M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module AO222M0HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO222M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module AO222M1HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO222M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module AO222M2HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO222M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module AO222M4HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO222M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module AO222M8HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO222M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B10M0HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B10M1HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B10M2HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B10M4HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B10M8HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B11M0HM_func( Z, A1, B1, NA2, NB2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, NA2, NB2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB2_org, NB2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B11M0HM_udp_0(Z,A1_org,NA2_org,B1_org,NB2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B11M1HM_func( Z, A1, B1, NA2, NB2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, NA2, NB2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB2_org, NB2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B11M0HM_udp_0(Z,A1_org,NA2_org,B1_org,NB2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B11M2HM_func( Z, A1, B1, NA2, NB2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, NA2, NB2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB2_org, NB2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B11M0HM_udp_0(Z,A1_org,NA2_org,B1_org,NB2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B11M4HM_func( Z, A1, B1, NA2, NB2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, NA2, NB2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB2_org, NB2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B11M0HM_udp_0(Z,A1_org,NA2_org,B1_org,NB2_org); 
endmodule
`endcelldefine

`celldefine
module AO22B11M8HM_func( Z, A1, B1, NA2, NB2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, NA2, NB2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB2_org, NB2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22B11M0HM_udp_0(Z,A1_org,NA2_org,B1_org,NB2_org); 
endmodule
`endcelldefine

`celldefine
module AO22M0HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22M1HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22M2HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22M4HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO22M8HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO31M0HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO31M1HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO31M1HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO31M1HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO31M2HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO31M1HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO31M4HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO31M1HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO31M8HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO31M1HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module AO32M0HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO32M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO32M1HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO32M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO32M2HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO32M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO32M4HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO32M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO32M8HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO32M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AO33M0HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO33M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module AO33M1HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO33M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module AO33M2HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO33M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module AO33M4HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO33M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module AO33M8HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AO33M1HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module AOI211M0HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI211M0HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI211M1HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI211M0HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI211M2HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI211M0HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI211M4HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI211M0HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI211M8HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI211M0HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B01M0HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B01M0HM_udp_0(Z,A1_org,NB_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B01M1HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B01M0HM_udp_0(Z,A1_org,NB_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B01M2HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B01M0HM_udp_0(Z,A1_org,NB_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B01M4HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B01M0HM_udp_0(Z,A1_org,NB_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B01M8HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B01M0HM_udp_0(Z,A1_org,NB_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B10M0HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B10M0HM_udp_0(Z,A1_org,B_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B10M1HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B10M0HM_udp_0(Z,A1_org,B_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B10M2HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B10M0HM_udp_0(Z,A1_org,B_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B10M4HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B10M0HM_udp_0(Z,A1_org,B_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B10M8HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B10M0HM_udp_0(Z,A1_org,B_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B20M0HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B20M1HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B20M2HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B20M4HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21B20M8HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M0HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M1HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M2HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M3HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M4HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M6HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI21M8HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI221M0HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI221M0HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI221M1HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI221M0HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI221M2HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI221M0HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI221M4HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI221M0HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI221M8HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI221M0HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI222M0HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI222M0HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI222M1HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI222M0HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI222M2HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI222M0HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI222M4HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI222M0HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI222M8HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI222M0HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22B20M0HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,B1_org,NA1_org,NA2_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22B20M1HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,B1_org,NA1_org,NA2_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22B20M2HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,B1_org,NA1_org,NA2_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22B20M4HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,B1_org,NA1_org,NA2_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22B20M8HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,B1_org,NA1_org,NA2_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22M0HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22M1HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22M2HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22M4HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI22M8HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module AOI31M0HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI31M0HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI31M1HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI31M0HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI31M2HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI31M0HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI31M4HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI31M0HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI31M8HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI31M0HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI32M0HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI32M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI32M1HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI32M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI32M2HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI32M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI32M4HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI32M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI32M8HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI32M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI33M0HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI33M0HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI33M1HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI33M0HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI33M2HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI33M0HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI33M4HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI33M0HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module AOI33M8HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI33M0HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module BUFM10HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM12HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM14HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM16HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM18HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM20HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM24HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM28HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM2HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM32HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM36HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM3HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM40HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM48HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM5HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM6HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFM8HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module BUFTM12HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM16HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM1HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM20HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM24HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM2HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM3HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM4HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM6HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module BUFTM8HM_func( Z, A, E, VDD , VSS );
inout VSS;
inout VDD;
input A, E;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0HM_udp_0(MGM_WB_0,A_org,E_org); 

	not MGM_BG_0(MGM_WB_1,E_org);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine

`celldefine
module CKAN2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKAN2M16HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKAN2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKAN2M3HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKAN2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKAN2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKAN2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKBUFM12HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM16HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM20HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM24HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM2HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM32HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM3HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM40HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM48HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM6HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKBUFM8HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM12HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM16HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM20HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM24HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM2HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM32HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM3HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM40HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM48HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM6HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKINVM8HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module CKMUX2M12HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKMUX2M2HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKMUX2M3HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKMUX2M4HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKMUX2M6HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKMUX2M8HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKND2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKND2M16HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKND2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKND2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKND2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKND2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKXOR2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKXOR2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKXOR2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKXOR2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module CKXOR2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module DEL1M1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL1M4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL2M1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL2M4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL3M1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL3M4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL4M1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DEL4M4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	buf MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module DFCM1HM_func( Q, QB, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCM2HM_func( Q, QB, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCM4HM_func( Q, QB, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCM8HM_func( Q, QB, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCQM1HM_func( Q, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQM2HM_func( Q, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQM4HM_func( Q, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQM8HM_func( Q, CKB, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQRSM1HM_func( Q, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQRSM2HM_func( Q, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQRSM4HM_func( Q, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCQRSM8HM_func( Q, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFCRSM1HM_func( Q, QB, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCRSM2HM_func( Q, QB, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCRSM4HM_func( Q, QB, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFCRSM8HM_func( Q, QB, CKB, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEM1HM_func( Q, QB, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEM2HM_func( Q, QB, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEM4HM_func( Q, QB, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEM8HM_func( Q, QB, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEQM1HM_func( Q, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQM2HM_func( Q, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQM4HM_func( Q, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQM8HM_func( Q, CK, D, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQRM1HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQRM2HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQRM4HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQRM8HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQZRM1HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQZRM2HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQZRM4HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFEQZRM8HM_func( Q, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFERM1HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFERM2HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFERM4HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFERM8HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	DFEM1HM_udp_0(MGM_D,D_org,E_org,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEZRM1HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEZRM2HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEZRM4HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFEZRM8HM_func( Q, QB, CK, D, E, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFM1HM_func( Q, QB, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFM2HM_func( Q, QB, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFM4HM_func( Q, QB, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFM8HM_func( Q, QB, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFMM1HM_func( Q, QB, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFMM2HM_func( Q, QB, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFMM4HM_func( Q, QB, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFMM8HM_func( Q, QB, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFMQM1HM_func( Q, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFMQM2HM_func( Q, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFMQM4HM_func( Q, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFMQM8HM_func( Q, CK, D1, D2, S,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	DFMM1HM_udp_0(MGM_D,D1_org,S_org,D2_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQM1HM_func( Q, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQM2HM_func( Q, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQM4HM_func( Q, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQM8HM_func( Q, CK, D,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRM1HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRM2HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRM4HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRM8HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRSM1HM_func( Q, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRSM2HM_func( Q, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRSM4HM_func( Q, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQRSM8HM_func( Q, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQSM1HM_func( Q, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQSM2HM_func( Q, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQSM4HM_func( Q, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQSM8HM_func( Q, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQZRM1HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQZRM2HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQZRM4HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFQZRM8HM_func( Q, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module DFRM1HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRM2HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRM4HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRM8HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRSM1HM_func( Q, QB, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRSM2HM_func( Q, QB, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRSM4HM_func( Q, QB, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFRSM8HM_func( Q, QB, CK, D, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,D_org,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFSM1HM_func( Q, QB, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFSM2HM_func( Q, QB, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFSM4HM_func( Q, QB, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFSM8HM_func( Q, QB, CK, D, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,D_org,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFZRM1HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFZRM2HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFZRM4HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module DFZRM8HM_func( Q, QB, CK, D, RB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_0(MGM_D,D_org,RB_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module INVM0HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM10HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM12HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM14HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM16HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM18HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM1HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM20HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM24HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM28HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM2HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM32HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM36HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM3HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM40HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM48HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM4HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM5HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM6HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module INVM8HM_func( Z, A, VDD , VSS );
inout VSS;
inout VDD;
input A;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(Z,A_org);
endmodule
`endcelldefine

`celldefine
module LACM0HM_func( Q, QB, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACM1HM_func( Q, QB, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACM2HM_func( Q, QB, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACM4HM_func( Q, QB, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACQM0HM_func( Q, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQM1HM_func( Q, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQM2HM_func( Q, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQM4HM_func( Q, D, GB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D_org,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQRSM0HM_func( Q, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQRSM1HM_func( Q, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQRSM2HM_func( Q, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACQRSM4HM_func( Q, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LACRSM0HM_func( Q, QB, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACRSM1HM_func( Q, QB, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACRSM2HM_func( Q, QB, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LACRSM4HM_func( Q, QB, D, GB, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, GB, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (GB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (GB_org, GB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_EN,GB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D_org,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LAGCECSM12HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL); 

endmodule
`endcelldefine

`celldefine
module LAGCECSM16HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL); 
 
endmodule
`endcelldefine

`celldefine
module LAGCECSM20HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL);
 
endmodule
`endcelldefine

`celldefine
module LAGCECSM2HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL);
 
endmodule
`endcelldefine

`celldefine
module LAGCECSM3HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL);
 
endmodule
`endcelldefine

`celldefine
module LAGCECSM4HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL); 
 
endmodule
`endcelldefine

`celldefine
module LAGCECSM6HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL);
 
endmodule
`endcelldefine

`celldefine
module LAGCECSM8HM_func( GCK, CKB, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, E, SE;
output GCK;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB_org,MGM_EN,notifier);
        not NGN_n0 (NOT_ENL, ENL);
	OR2M0HM_udp_0(GCK,CKB_org,NOT_ENL);
 
endmodule
`endcelldefine

`celldefine
module LAGCEM12HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM16HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM20HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM2HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM3HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM4HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM6HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCEM8HM_func( GCK, CK, E,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,E_org,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM12HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM16HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM20HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM2HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM3HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM4HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM6HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAGCESM8HM_func( GCK, CK, E, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, E, SE;
output GCK;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));
 
        OR2M0HM_udp_0(MGM_EN,E_org,SE_org); 
        not NGN_n0 (CKB, CK_org);
        MGM_IQ_LATCH_UDP(ENL,1'b0,1'b0,CKB,MGM_EN,notifier);
	ADHM1HM_udp_0(GCK,CK_org,ENL); 
endmodule
`endcelldefine

`celldefine
module LAM0HM_func( Q, QB, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LAM1HM_func( Q, QB, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LAM2HM_func( Q, QB, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LAM4HM_func( Q, QB, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LAQM0HM_func( Q, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQM1HM_func( Q, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQM2HM_func( Q, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQM4HM_func( Q, D, G,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G_org,D_org,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G_org,D_org,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQRSM0HM_func( Q, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQRSM1HM_func( Q, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQRSM2HM_func( Q, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LAQRSM4HM_func( Q, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module LARSM0HM_func( Q, QB, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LARSM1HM_func( Q, QB, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LARSM2HM_func( Q, QB, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module LARSM4HM_func( Q, QB, D, G, RB, SB,notifier, VDD , VSS );
inout VSS;
inout VDD;
input D, G, RB, SB;
output Q, QB;
input notifier;
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (G_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (G_org, G, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G_org,D_org,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G_org,D_org,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module MAO222M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAO222M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAO222M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAO222M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AD42M2HM_udp_1(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAOI2223M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MAOI2223M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MAOI2223M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MAOI2223M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MAOI2223M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MAOI2223M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MAOI2223M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MAOI2223M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MAOI222M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAOI222M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAOI222M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAOI222M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MAOI22M0HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module MAOI22M1HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module MAOI22M2HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module MAOI22M4HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	AOI22B20M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module MOAI22M0HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module MOAI22M1HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module MOAI22M2HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module MOAI22M4HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M0HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M1HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M2HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M3HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M4HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M6HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX2M8HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MUX3M0HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MUX3M1HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MUX3M2HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MUX3M4HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MUX4M0HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MUX4M1HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MUX4M2HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MUX4M4HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MUX4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M0HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M1HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M2HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M3HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M4HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M6HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB2M8HM_func( Z, A, B, S, VDD , VSS );
inout VSS;
inout VDD;
input A, B, S;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB2M0HM_udp_0(Z,A_org,S_org,B_org); 
endmodule
`endcelldefine

`celldefine
module MXB3M0HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MXB3M1HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MXB3M2HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MXB3M4HM_func( Z, A, B, C, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB3M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module MXB4M0HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MXB4M1HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MXB4M2HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module MXB4M4HM_func( Z, A, B, C, D, S0, S1, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, S0, S1;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S0_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S0_org, S0, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S1_org, S1, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MXB4M0HM_udp_0(Z,A_org,S0_org,S1_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND2B1M0HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND2B1M12HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND2B1M1HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND2B1M2HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND2B1M4HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND2B1M8HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND2M0HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M16HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M3HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M5HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module ND3B1M0HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND3B1M1HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND3B1M2HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND3B1M4HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND3B1M8HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND3M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M12HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M16HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M3HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M6HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND3M8HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module ND4B1M0HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND4B1M1HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND4B1M2HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND4B1M4HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND4B1M8HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module ND4B2M0HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module ND4B2M1HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module ND4B2M2HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module ND4B2M4HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module ND4B2M8HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module ND4M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M12HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M16HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M6HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module ND4M8HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ND4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR2B1M0HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR2B1M12HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR2B1M1HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR2B1M2HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR2B1M4HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR2B1M8HM_func( Z, B, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR2B1M0HM_udp_0(Z,B_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR2M0HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M16HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M3HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M5HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADCSIOM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module NR3B1M0HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR3B1M1HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR3B1M2HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR3B1M4HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR3B1M8HM_func( Z, B, C, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3B1M0HM_udp_0(Z,B_org,C_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR3M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M12HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M16HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M6HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR3M8HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module NR4B1M0HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR4B1M1HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR4B1M2HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR4B1M4HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR4B1M8HM_func( Z, B, C, D, NA, VDD , VSS );
inout VSS;
inout VDD;
input B, C, D, NA;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B1M0HM_udp_0(Z,B_org,C_org,D_org,NA_org); 
endmodule
`endcelldefine

`celldefine
module NR4B2M0HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module NR4B2M1HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module NR4B2M2HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module NR4B2M4HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module NR4B2M8HM_func( Z, C, D, NA, NB, VDD , VSS );
inout VSS;
inout VDD;
input C, D, NA, NB;
output Z;
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA_org, NA, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4B2M0HM_udp_0(Z,C_org,D_org,NA_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module NR4M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M12HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M16HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M6HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module NR4M8HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	NR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OA211M0HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA211M12HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA211M1HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA211M12HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA211M2HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA211M12HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA211M4HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA211M12HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA211M8HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA211M12HM_udp_0(Z,A1_org,B_org,C_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA21M0HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA21M1HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA21M2HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA21M4HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA21M8HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA21M0HM_udp_0(Z,A1_org,B_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA221M0HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA221M1HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA221M1HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA221M1HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA221M2HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA221M1HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA221M4HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA221M1HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA221M8HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA221M1HM_udp_0(Z,A1_org,B1_org,C_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA222M0HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA222M1HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA222M1HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA222M1HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA222M2HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA222M1HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA222M4HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA222M1HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA222M8HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA222M1HM_udp_0(Z,A1_org,B1_org,C1_org,C2_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA22M0HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA22M1HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA22M2HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA22M4HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA22M8HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA22M0HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org); 
endmodule
`endcelldefine

`celldefine
module OA31M0HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA31M1HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA31M1HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA31M1HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA31M2HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA31M1HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA31M4HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA31M1HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA31M8HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA31M1HM_udp_0(Z,A1_org,B_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA32M0HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA32M1HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA32M1HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA32M1HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA32M2HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA32M1HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA32M4HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA32M1HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA32M8HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA32M1HM_udp_0(Z,A1_org,B1_org,B2_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA33M0HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA33M1HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA33M1HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA33M1HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA33M2HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA33M1HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA33M4HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA33M1HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OA33M8HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OA33M1HM_udp_0(Z,A1_org,B1_org,B2_org,B3_org,A2_org,A3_org); 
endmodule
`endcelldefine

`celldefine
module OAI211B100M0HM_func( Z, A1, B, C, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, C, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211B100M0HM_udp_0(Z,A1_org,NA2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211B100M1HM_func( Z, A1, B, C, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, C, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211B100M0HM_udp_0(Z,A1_org,NA2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211B100M2HM_func( Z, A1, B, C, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, C, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211B100M0HM_udp_0(Z,A1_org,NA2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211B100M4HM_func( Z, A1, B, C, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, C, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211B100M0HM_udp_0(Z,A1_org,NA2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211B100M8HM_func( Z, A1, B, C, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, C, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211B100M0HM_udp_0(Z,A1_org,NA2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211M0HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211M0HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211M1HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211M0HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211M2HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211M0HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211M4HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211M0HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI211M8HM_func( Z, A1, A2, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI211M0HM_udp_0(Z,A1_org,A2_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B01M0HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	BEM2HM_udp_1(Z,A1_org,A2_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B01M1HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	BEM2HM_udp_1(Z,A1_org,A2_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B01M2HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	BEM2HM_udp_1(Z,A1_org,A2_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B01M4HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	BEM2HM_udp_1(Z,A1_org,A2_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B01M8HM_func( Z, A1, A2, NB, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, NB;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NB_org, NB, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	BEM2HM_udp_1(Z,A1_org,A2_org,NB_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B10M0HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B10M0HM_udp_0(Z,A1_org,NA2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B10M1HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B10M0HM_udp_0(Z,A1_org,NA2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B10M2HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B10M0HM_udp_0(Z,A1_org,NA2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B10M4HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B10M0HM_udp_0(Z,A1_org,NA2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B10M8HM_func( Z, A1, B, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B10M0HM_udp_0(Z,A1_org,NA2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B20M0HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B20M1HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B20M2HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B20M4HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI21B20M8HM_func( Z, B, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B, NA1, NA2;
output Z;
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21B20M0HM_udp_0(Z,B_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M0HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M1HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M2HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M3HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M4HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M6HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI21M8HM_func( Z, A1, A2, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI21M0HM_udp_0(Z,A1_org,A2_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI221M0HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI221M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI221M1HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI221M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI221M2HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI221M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI221M4HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI221M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI221M8HM_func( Z, A1, A2, B1, B2, C, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI221M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OAI222M0HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI222M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module OAI222M1HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI222M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module OAI222M2HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI222M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module OAI222M4HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI222M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module OAI222M8HM_func( Z, A1, A2, B1, B2, C1, C2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2, C1, C2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C1_org, C1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C2_org, C2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI222M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org,C1_org,C2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B10M0HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B10M1HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B10M2HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B10M4HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B10M8HM_func( Z, A1, B1, B2, NA2, VDD , VSS );
inout VSS;
inout VDD;
input A1, B1, B2, NA2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22B10M0HM_udp_0(Z,A1_org,NA2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B20M0HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,B1_org,B2_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B20M1HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,B1_org,B2_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B20M2HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,B1_org,B2_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B20M4HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,B1_org,B2_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22B20M8HM_func( Z, B1, B2, NA1, NA2, VDD , VSS );
inout VSS;
inout VDD;
input B1, B2, NA1, NA2;
output Z;
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA1_org, NA1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (NA2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (NA2_org, NA2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	MOAI22M1HM_udp_0(Z,B1_org,B2_org,NA1_org,NA2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22M0HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22M1HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22M2HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22M4HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI22M8HM_func( Z, A1, A2, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI22M0HM_udp_0(Z,A1_org,A2_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI31M0HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI31M0HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI31M1HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI31M0HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI31M2HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI31M0HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI31M4HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI31M0HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI31M8HM_func( Z, A1, A2, A3, B, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI31M0HM_udp_0(Z,A1_org,A2_org,A3_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OAI32M0HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI32M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI32M1HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI32M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI32M2HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI32M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI32M4HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI32M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI32M8HM_func( Z, A1, A2, A3, B1, B2, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI32M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org); 
endmodule
`endcelldefine

`celldefine
module OAI33M0HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI33M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module OAI33M1HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI33M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module OAI33M2HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI33M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module OAI33M4HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI33M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module OAI33M8HM_func( Z, A1, A2, A3, B1, B2, B3, VDD , VSS );
inout VSS;
inout VDD;
input A1, A2, A3, B1, B2, B3;
output Z;
bufif1 (A1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A1_org, A1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A2_org, A2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (A3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A3_org, A3, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B1_org, B1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B2_org, B2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B3_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B3_org, B3, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OAI33M0HM_udp_0(Z,A1_org,A2_org,A3_org,B1_org,B2_org,B3_org); 
endmodule
`endcelldefine

`celldefine
module OR2M0HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M12HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M16HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR2M0HM_udp_0(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module OR3M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M12HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M16HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M6HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR3M8HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR3M0HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module OR4M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M12HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M16HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M6HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR4M8HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR4M0HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module OR6M0HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module OR6M12HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module OR6M1HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module OR6M2HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module OR6M4HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module OR6M6HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module OR6M8HM_func( Z, A, B, C, D, E, F, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D, E, F;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (F_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (F_org, F, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	OR6M12HM_udp_0(Z,A_org,B_org,C_org,D_org,E_org,F_org); 
endmodule
`endcelldefine

`celldefine
module SDFCM1HM_func( Q, QB, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCM2HM_func( Q, QB, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCM4HM_func( Q, QB, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCM8HM_func( Q, QB, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCQM1HM_func( Q, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQM2HM_func( Q, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQM4HM_func( Q, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQM8HM_func( Q, CKB, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQRSM1HM_func( Q, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQRSM2HM_func( Q, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQRSM4HM_func( Q, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCQRSM8HM_func( Q, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFCRSM1HM_func( Q, QB, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCRSM2HM_func( Q, QB, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCRSM4HM_func( Q, QB, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFCRSM8HM_func( Q, QB, CKB, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CKB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CKB_org, CKB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_CLK,CKB_org);

	not MGM_BG_1(MGM_P,SB_org);

	not MGM_BG_2(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEM1HM_func( Q, QB, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEM2HM_func( Q, QB, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEM4HM_func( Q, QB, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEM8HM_func( Q, QB, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEQM1HM_func( Q, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQM2HM_func( Q, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQM4HM_func( Q, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQM8HM_func( Q, CK, D, E, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQRM1HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQRM2HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQRM4HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQRM8HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQZRM1HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQZRM2HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQZRM4HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFEQZRM8HM_func( Q, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFERM1HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFERM2HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFERM4HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFERM8HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	SDFEM1HM_udp_0(MGM_D,D_org,E_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEZRM1HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEZRM2HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEZRM4HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFEZRM8HM_func( Q, QB, CK, D, E, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (E_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (E_org, E, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFEQZRM1HM_udp_0(MGM_D,D_org,E_org,RB_org,SE_org,IQ,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFM1HM_func( Q, QB, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFM2HM_func( Q, QB, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFM4HM_func( Q, QB, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFM8HM_func( Q, QB, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFMM1HM_func( Q, QB, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFMM2HM_func( Q, QB, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFMM4HM_func( Q, QB, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFMM8HM_func( Q, QB, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFMQM1HM_func( Q, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFMQM2HM_func( Q, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFMQM4HM_func( Q, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFMQM8HM_func( Q, CK, D1, D2, S, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D1_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D1_org, D1, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D2_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D2_org, D2, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (S_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (S_org, S, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFMM1HM_udp_0(MGM_D,D1_org,S_org,SE_org,D2_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQM1HM_func( Q, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQM2HM_func( Q, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQM4HM_func( Q, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQM8HM_func( Q, CK, D, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRM1HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRM2HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRM4HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRM8HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRSM1HM_func( Q, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRSM2HM_func( Q, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRSM4HM_func( Q, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRSM8HM_func( Q, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQRXM2HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQSM1HM_func( Q, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQSM2HM_func( Q, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQSM4HM_func( Q, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQSM8HM_func( Q, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQZRM1HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQZRM2HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQZRM4HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFQZRM8HM_func( Q, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine

`celldefine
module SDFRM1HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRM2HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRM4HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRM8HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRSM1HM_func( Q, QB, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRSM2HM_func( Q, QB, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRSM4HM_func( Q, QB, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFRSM8HM_func( Q, QB, CK, D, RB, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	not MGM_BG_1(MGM_C,RB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFSM1HM_func( Q, QB, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFSM2HM_func( Q, QB, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFSM4HM_func( Q, QB, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFSM8HM_func( Q, QB, CK, D, SB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SB_org, SB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	not MGM_BG_0(MGM_P,SB_org);

	CKMUX2M12HM_udp_0(MGM_D,D_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK_org,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFZRM1HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFZRM2HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFZRM4HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module SDFZRM8HM_func( Q, QB, CK, D, RB, SD, SE,notifier, VDD , VSS );
inout VSS;
inout VDD;
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;
bufif1 (CK_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (CK_org, CK, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (RB_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (RB_org, RB, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SD_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SD_org, SD, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (SE_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (SE_org, SE, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	SDFAQM1HM_udp_0(MGM_D,D_org,RB_org,SE_org,SD_org); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK_org,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK_org,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine

`celldefine
module TIE0HM_func( Z, VDD , VSS );
inout VSS;
inout VDD;
output Z;

        buf I0 (out_temp, 1'b0);
	assign Z = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

endmodule
`endcelldefine

`celldefine
module TIE1HM_func( Z, VDD , VSS );
inout VSS;
inout VDD;
output Z;

        buf I1 (out_temp, 1'b1);
	assign Z = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;	
endmodule
`endcelldefine

`celldefine
module XNR2M0HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHCM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XNR2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHCM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XNR2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHCM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XNR2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHCM2HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XNR3M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XNR3M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XNR3M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XNR3M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XNR4M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XNR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XNR4M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XNR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XNR4M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XNR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XNR4M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XNR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M0HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M1HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M2HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M3HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M4HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M6HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR2M8HM_func( Z, A, B, VDD , VSS );
inout VSS;
inout VDD;
input A, B;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADHM1HM_udp_1(Z,A_org,B_org); 
endmodule
`endcelldefine

`celldefine
module XOR3M0HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCSIOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XOR3M1HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCSIOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XOR3M2HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCSIOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XOR3M4HM_func( Z, A, B, C, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	ADFCSIOM2HM_udp_0(Z,A_org,B_org,C_org); 
endmodule
`endcelldefine

`celldefine
module XOR4M0HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XOR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XOR4M1HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XOR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XOR4M2HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XOR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine

`celldefine
module XOR4M4HM_func( Z, A, B, C, D, VDD , VSS );
inout VSS;
inout VDD;
input A, B, C, D;
output Z;
bufif1 (A_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (A_org, A, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (B_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (B_org, B, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (C_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (C_org, C, ((VDD !== 1'b1) || (VSS !== 1'b0)));
bufif1 (D_org, 1'bx, ((VDD !== 1'b1) || (VSS !== 1'b0) ));
bufif0 (D_org, D, ((VDD !== 1'b1) || (VSS !== 1'b0)));

	XOR4M1HM_udp_0(Z,A_org,B_org,C_org,D_org); 
endmodule
`endcelldefine


primitive AD42M2HM_udp_1(ICO,A, B, C);
  output ICO;
  input A, B, C;
  table
  //A, B, C: ICO
    1  1  ?: 1;
    1  ?  1: 1;
    ?  1  1: 1;
    0  0  ?: 0;
    0  ?  0: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive ADCSIOM2HM_udp_0(CO0B,A, B);
  output CO0B;
  input A, B;
  table
  //A, B: CO0B
    0  ?: 1;
    ?  0: 1;
    1  1: 0;
  endtable
endprimitive

primitive ADCSIOM2HM_udp_1(CO1B,A, B);
  output CO1B;
  input A, B;
  table
  //A, B: CO1B
    0  0: 1;
    1  ?: 0;
    ?  1: 0;
  endtable
endprimitive

primitive ADCSOM2HM_udp_0(CO0B,A, B, CI0);
  output CO0B;
  input A, B, CI0;
  table
  //A, B, CI0: CO0B
    0  0  ?: 1;
    0  ?  0: 1;
    ?  0  0: 1;
    1  1  ?: 0;
    1  ?  1: 0;
    ?  1  1: 0;
  endtable
endprimitive

primitive ADFCM2HM_udp_0(S,A, B, NCI);
  output S;
  input A, B, NCI;
  table
  //A, B, NCI: S
    1  1  0: 1;
    1  0  1: 1;
    0  1  1: 1;
    0  0  0: 1;
    1  1  1: 0;
    1  0  0: 0;
    0  1  0: 0;
    0  0  1: 0;
  endtable
endprimitive

primitive ADFCSIOM2HM_udp_0(S,A, B, CS);
  output S;
  input A, B, CS;
  table
  //A, B, CS: S
    1  1  1: 1;
    1  0  0: 1;
    0  1  0: 1;
    0  0  1: 1;
    1  1  0: 0;
    1  0  1: 0;
    0  1  1: 0;
    0  0  0: 0;
  endtable
endprimitive

primitive ADHCM2HM_udp_1(S,A, NCI);
  output S;
  input A, NCI;
  table
  //A, NCI: S
    1  1: 1;
    0  0: 1;
    1  0: 0;
    0  1: 0;
  endtable
endprimitive

primitive ADHM1HM_udp_0(CO,A, B);
  output CO;
  input A, B;
  table
  //A, B: CO
    1  1: 1;
    0  ?: 0;
    ?  0: 0;
  endtable
endprimitive

primitive ADHM1HM_udp_1(S,A, B);
  output S;
  input A, B;
  table
  //A, B: S
    1  0: 1;
    0  1: 1;
    1  1: 0;
    0  0: 0;
  endtable
endprimitive

primitive AN3M0HM_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    1  1  1: 1;
    0  ?  ?: 0;
    ?  0  ?: 0;
    ?  ?  0: 0;
  endtable
endprimitive

primitive AN4M0HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  1  1  1: 1;
    0  ?  ?  ?: 0;
    ?  0  ?  ?: 0;
    ?  ?  0  ?: 0;
    ?  ?  ?  0: 0;
  endtable
endprimitive

primitive AO211M1HM_udp_0(Z,A1, A2, B, C);
  output Z;
  input A1, A2, B, C;
  table
  //A1, A2, B, C: Z
    1  1  ?  ?: 1;
    ?  ?  1  ?: 1;
    ?  ?  ?  1: 1;
    0  ?  0  0: 0;
    ?  0  0  0: 0;
  endtable
endprimitive

primitive AO21M0HM_udp_0(Z,A1, A2, B);
  output Z;
  input A1, A2, B;
  table
  //A1, A2, B: Z
    1  1  ?: 1;
    ?  ?  1: 1;
    0  ?  0: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive AO221M1HM_udp_0(Z,A1, A2, B1, B2, C);
  output Z;
  input A1, A2, B1, B2, C;
  table
  //A1, A2, B1, B2, C: Z
    1  1  ?  ?  ?: 1;
    ?  ?  1  1  ?: 1;
    ?  ?  ?  ?  1: 1;
    0  ?  0  ?  0: 0;
    0  ?  ?  0  0: 0;
    ?  0  0  ?  0: 0;
    ?  0  ?  0  0: 0;
  endtable
endprimitive

primitive AO222M1HM_udp_0(Z,A1, A2, B1, B2, C1, C2);
  output Z;
  input A1, A2, B1, B2, C1, C2;
  table
  //A1, A2, B1, B2, C1, C2: Z
    1  1  ?  ?  ?  ?: 1;
    ?  ?  1  1  ?  ?: 1;
    ?  ?  ?  ?  1  1: 1;
    0  ?  0  ?  0  ?: 0;
    0  ?  0  ?  ?  0: 0;
    0  ?  ?  0  0  ?: 0;
    0  ?  ?  0  ?  0: 0;
    ?  0  0  ?  0  ?: 0;
    ?  0  0  ?  ?  0: 0;
    ?  0  ?  0  0  ?: 0;
    ?  0  ?  0  ?  0: 0;
  endtable
endprimitive

primitive AO22B10M0HM_udp_0(Z,A1, NA2, B1, B2);
  output Z;
  input A1, NA2, B1, B2;
  table
  //A1, NA2, B1, B2: Z
    1  0  ?  ?: 1;
    ?  ?  1  1: 1;
    0  ?  0  ?: 0;
    0  ?  ?  0: 0;
    ?  1  0  ?: 0;
    ?  1  ?  0: 0;
  endtable
endprimitive

primitive AO22B11M0HM_udp_0(Z,A1, NA2, B1, NB2);
  output Z;
  input A1, NA2, B1, NB2;
  table
  //A1, NA2, B1, NB2: Z
    1  0  ?  ?: 1;
    ?  ?  1  0: 1;
    0  ?  0  ?: 0;
    0  ?  ?  1: 0;
    ?  1  0  ?: 0;
    ?  1  ?  1: 0;
  endtable
endprimitive

primitive AO22M0HM_udp_0(Z,A1, A2, B1, B2);
  output Z;
  input A1, A2, B1, B2;
  table
  //A1, A2, B1, B2: Z
    1  1  ?  ?: 1;
    ?  ?  1  1: 1;
    0  ?  0  ?: 0;
    0  ?  ?  0: 0;
    ?  0  0  ?: 0;
    ?  0  ?  0: 0;
  endtable
endprimitive

primitive AO31M1HM_udp_0(Z,A1, A2, A3, B);
  output Z;
  input A1, A2, A3, B;
  table
  //A1, A2, A3, B: Z
    1  1  1  ?: 1;
    ?  ?  ?  1: 1;
    0  ?  ?  0: 0;
    ?  0  ?  0: 0;
    ?  ?  0  0: 0;
  endtable
endprimitive

primitive AO32M1HM_udp_0(Z,A1, A2, A3, B1, B2);
  output Z;
  input A1, A2, A3, B1, B2;
  table
  //A1, A2, A3, B1, B2: Z
    1  1  1  ?  ?: 1;
    ?  ?  ?  1  1: 1;
    0  ?  ?  0  ?: 0;
    0  ?  ?  ?  0: 0;
    ?  0  ?  0  ?: 0;
    ?  0  ?  ?  0: 0;
    ?  ?  0  0  ?: 0;
    ?  ?  0  ?  0: 0;
  endtable
endprimitive

primitive AO33M1HM_udp_0(Z,A1, A2, A3, B1, B2, B3);
  output Z;
  input A1, A2, A3, B1, B2, B3;
  table
  //A1, A2, A3, B1, B2, B3: Z
    1  1  1  ?  ?  ?: 1;
    ?  ?  ?  1  1  1: 1;
    0  ?  ?  0  ?  ?: 0;
    0  ?  ?  ?  0  ?: 0;
    0  ?  ?  ?  ?  0: 0;
    ?  0  ?  0  ?  ?: 0;
    ?  0  ?  ?  0  ?: 0;
    ?  0  ?  ?  ?  0: 0;
    ?  ?  0  0  ?  ?: 0;
    ?  ?  0  ?  0  ?: 0;
    ?  ?  0  ?  ?  0: 0;
  endtable
endprimitive

primitive AOI211M0HM_udp_0(Z,A1, B, C, A2);
  output Z;
  input A1, B, C, A2;
  table
  //A1, B, C, A2: Z
    0  0  0  ?: 1;
    ?  0  0  0: 1;
    1  ?  ?  1: 0;
    ?  1  ?  ?: 0;
    ?  ?  1  ?: 0;
  endtable
endprimitive

primitive AOI21B01M0HM_udp_0(Z,A1, NB, A2);
  output Z;
  input A1, NB, A2;
  table
  //A1, NB, A2: Z
    0  1  ?: 1;
    ?  1  0: 1;
    1  ?  1: 0;
    ?  0  ?: 0;
  endtable
endprimitive

primitive AOI21B10M0HM_udp_0(Z,A1, B, NA2);
  output Z;
  input A1, B, NA2;
  table
  //A1, B, NA2: Z
    0  0  ?: 1;
    ?  0  1: 1;
    1  ?  0: 0;
    ?  1  ?: 0;
  endtable
endprimitive

primitive AOI21B20M0HM_udp_0(Z,B, NA1, NA2);
  output Z;
  input B, NA1, NA2;
  table
  //B, NA1, NA2: Z
    0  1  ?: 1;
    0  ?  1: 1;
    1  ?  ?: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive AOI21M0HM_udp_0(Z,A1, B, A2);
  output Z;
  input A1, B, A2;
  table
  //A1, B, A2: Z
    0  0  ?: 1;
    ?  0  0: 1;
    1  ?  1: 0;
    ?  1  ?: 0;
  endtable
endprimitive

primitive AOI221M0HM_udp_0(Z,A1, B1, C, B2, A2);
  output Z;
  input A1, B1, C, B2, A2;
  table
  //A1, B1, C, B2, A2: Z
    0  0  0  ?  ?: 1;
    0  ?  0  0  ?: 1;
    ?  0  0  ?  0: 1;
    ?  ?  0  0  0: 1;
    1  ?  ?  ?  1: 0;
    ?  1  ?  1  ?: 0;
    ?  ?  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI222M0HM_udp_0(Z,A1, B1, C1, C2, B2, A2);
  output Z;
  input A1, B1, C1, C2, B2, A2;
  table
  //A1, B1, C1, C2, B2, A2: Z
    0  0  0  ?  ?  ?: 1;
    0  0  ?  0  ?  ?: 1;
    0  ?  0  ?  0  ?: 1;
    0  ?  ?  0  0  ?: 1;
    ?  0  0  ?  ?  0: 1;
    ?  0  ?  0  ?  0: 1;
    ?  ?  0  ?  0  0: 1;
    ?  ?  ?  0  0  0: 1;
    1  ?  ?  ?  ?  1: 0;
    ?  1  ?  ?  1  ?: 0;
    ?  ?  1  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI22B20M0HM_udp_0(Z,B1, NA1, NA2, B2);
  output Z;
  input B1, NA1, NA2, B2;
  table
  //B1, NA1, NA2, B2: Z
    0  1  ?  ?: 1;
    0  ?  1  ?: 1;
    ?  1  ?  0: 1;
    ?  ?  1  0: 1;
    1  ?  ?  1: 0;
    ?  0  0  ?: 0;
  endtable
endprimitive

primitive AOI22M0HM_udp_0(Z,A1, B1, B2, A2);
  output Z;
  input A1, B1, B2, A2;
  table
  //A1, B1, B2, A2: Z
    0  0  ?  ?: 1;
    0  ?  0  ?: 1;
    ?  0  ?  0: 1;
    ?  ?  0  0: 1;
    1  ?  ?  1: 0;
    ?  1  1  ?: 0;
  endtable
endprimitive

primitive AOI31M0HM_udp_0(Z,A1, B, A2, A3);
  output Z;
  input A1, B, A2, A3;
  table
  //A1, B, A2, A3: Z
    0  0  ?  ?: 1;
    ?  0  0  ?: 1;
    ?  0  ?  0: 1;
    1  ?  1  1: 0;
    ?  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI32M0HM_udp_0(Z,A1, B1, B2, A2, A3);
  output Z;
  input A1, B1, B2, A2, A3;
  table
  //A1, B1, B2, A2, A3: Z
    0  0  ?  ?  ?: 1;
    0  ?  0  ?  ?: 1;
    ?  0  ?  0  ?: 1;
    ?  ?  0  0  ?: 1;
    ?  0  ?  ?  0: 1;
    ?  ?  0  ?  0: 1;
    1  ?  ?  1  1: 0;
    ?  1  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI33M0HM_udp_0(Z,A1, B1, B2, B3, A2, A3);
  output Z;
  input A1, B1, B2, B3, A2, A3;
  table
  //A1, B1, B2, B3, A2, A3: Z
    0  0  ?  ?  ?  ?: 1;
    0  ?  0  ?  ?  ?: 1;
    0  ?  ?  0  ?  ?: 1;
    ?  0  ?  ?  0  ?: 1;
    ?  ?  0  ?  0  ?: 1;
    ?  ?  ?  0  0  ?: 1;
    ?  0  ?  ?  ?  0: 1;
    ?  ?  0  ?  ?  0: 1;
    ?  ?  ?  0  ?  0: 1;
    1  ?  ?  ?  1  1: 0;
    ?  1  1  1  ?  ?: 0;
  endtable
endprimitive

primitive BEM2HM_udp_1(OA2,M0, M1, M2);
  output OA2;
  input M0, M1, M2;
  table
  //M0, M1, M2: OA2
    0  0  ?: 1;
    ?  ?  1: 1;
    1  ?  0: 0;
    ?  1  0: 0;
  endtable
endprimitive

primitive BUFTM0HM_udp_0(MGM_WB_0,A, E);
  output MGM_WB_0;
  input A, E;
  table
  //A, E: MGM_WB_0
    1  1: 1;
    0  1: 0;
    ?  0: 1;   
  endtable
endprimitive

primitive CKMUX2M12HM_udp_0(Z,A, S, B);
  output Z;
  input A, S, B;
  table
  //A, S, B: Z
    1  0  ?: 1;
    ?  1  1: 1;
    0  0  ?: 0;
    ?  1  0: 0;
    1  ?  1: 1;
    0  ?  0: 0;
  endtable
endprimitive

primitive DFEM1HM_udp_0(MGM_D,D, E, IQ);
  output MGM_D;
  input D, E, IQ;
  table
  //D, E, IQ: MGM_D
    1  1  ?: 1;
    1  ?  1: 1;
    ?  0  1: 1;
    0  1  ?: 0;
    0  ?  0: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive DFEQZRM1HM_udp_0(MGM_D,D, E, RB, IQ);
  output MGM_D;
  input D, E, RB, IQ;
  table
  //D, E, RB, IQ: MGM_D
    1  1  1  ?: 1;
    1  ?  1  1: 1;
    ?  0  1  1: 1;
    0  1  ?  ?: 0;
    0  ?  ?  0: 0;
    ?  0  ?  0: 0;
    ?  ?  0  ?: 0;
  endtable
endprimitive

primitive DFMM1HM_udp_0(MGM_D,D1, S, D2);
  output MGM_D;
  input D1, S, D2;
  table
  //D1, S, D2: MGM_D
    1  1  ?: 1;
    ?  0  1: 1;
    0  1  ?: 0;
    ?  0  0: 0;
    1  ?  1: 1;
    0  ?  0: 0;
  endtable
endprimitive

primitive MAOI2223M1HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    0  0  0  ?: 1;
    0  ?  ?  0: 1;
    ?  0  ?  0: 1;
    ?  ?  0  0: 1;
    1  1  1  ?: 0;
    1  ?  ?  1: 0;
    ?  1  ?  1: 0;
    ?  ?  1  1: 0;
  endtable
endprimitive

primitive MGM_H_IQ_LATCH_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  Q  :  Q 
  ?  ?  0  *  ?  :  ?  :  -;  // No change CK=0
  ?  0  1  0  ?  :  ?  :  0;  // Latch 0 
  ?  0  *  0  ?  :  0  :  0;  // reduce pessimism when D=0
  1  0  ?  ?  ?  :  ?  :  0;  // clear
  0  ?  1  1  ?  :  ?  :  1;  // Latch 1
  0  ?  *  1  ?  :  1  :  1;  // reduce pessimism when D=1
  ?  1  ?  ?  ?  :  ?  :  1;  // Preset P dominate C
  *  0  0  ?  ?  :  0  :  0;   // reduce clear pessimism
  *  0  ?  0  ?  :  0  :  0;   // reduce clear pessimism
  0  *  0  ?  ?  :  1  :  1;   // reduce preset pessimism
  0  *  ?  1  ?  :  1  :  1;   // reduce preset pessimism

//  ?  ?  ?  ?  *  :  ?  :  x;  // notifier
                  
endtable
endprimitive

primitive MGM_H_IQN_FF_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  QN  :  QN 
  ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  1;  // CK in 0
  ?  0  p  0  ?  :  1  :  1;  // reduce pessimism D=0
  1  ?  ?  ?  ?  :  ?  :  1;  // clear: C dominate P
  0  ?  r  1  ?  :  ?  :  0;  // CK in 1
  0  ?  p  1  ?  :  0  :  0;  // reduce pessimism D=1
  0  1  ?  ?  ?  :  ?  :  0;  // preset
  ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
  *  0  b  ?  ?  :  1  :  1;  // reduce clear pessimism
  *  0  x  0  ?  :  1  :  1;  // reduce clear pessimism
  0  *  b  ?  ?  :  0  :  0;  // reduce preset pessimism
  0  *  x  1  ?  :  0  :  0;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_IQ_FF_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//  C  P  CK  D  N :  Q  :  Q 
    ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
    ?  0  r  0  ?  :  ?  :  0;  // CK in 0
    ?  0  p  0  ?  :  0  :  0;  // reduce pessimism D=0
    1  ?  ?  ?  ?  :  ?  :  0;  // clear: C dominate P
    0  ?  r  1  ?  :  ?  :  1;  // CK in 1
    0  ?  p  1  ?  :  1  :  1;  // reduce pessimism D=1
    0  1  ?  ?  ?  :  ?  :  1;  // preset
    ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
    *  0  b  ?  ?  :  0  :  0;  // reduce clear pessimism
    *  0  x  0  ?  :  0  :  0;  // reduce clear pessimism
    0  *  b  ?  ?  :  1  :  1;  // reduce preset pessimism
    0  *  x  1  ?  :  1  :  1;  // reduce preset pessimism
//  ?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_IQ_LATCH_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//  C  P  CK  D  N :  Q  :  Q 
    ?  ?  0  *  ?  :  ?  :  -;   // No change CK=0
    ?  0  1  0  ?  :  ?  :  0;   // Latch 0
    ?  0  *  0  ?  :  0  :  0;   // reduce pessimism when D=0
    1  ?  ?  ?  ?  :  ?  :  0;   // Clear : C dominate P
    0  ?  1  1  ?  :  ?  :  1;   // Latch 1
    0  ?  *  1  ?  :  1  :  1;   // reduce pessimism when D=1
    0  1  ?  ?  ?  :  ?  :  1;   // Preset
    *  0  0  ?  ?  :  0  :  0;   // reduce clear pessimism
    *  0  ?  0  ?  :  0  :  0;   // reduce clear pessimism
    0  *  0  ?  ?  :  1  :  1;   // reduce preset pessimism
    0  *  ?  1  ?  :  1  :  1;   // reduce preset pessimism
//  ?  ?  ?  ?  *  :  ?  :  x;   // notifier
                  
endtable
endprimitive

primitive MGM_IQN_FF_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  QN  :  QN 
  ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  1;  // CK in 0
  ?  0  p  0  ?  :  1  :  1;  // reduce pessimism D=0
  1  ?  ?  ?  ?  :  ?  :  1;  // clear: C dominate P
  0  ?  r  1  ?  :  ?  :  0;  // CK in 1
  0  ?  p  1  ?  :  0  :  0;  // reduce pessimism D=1
  0  1  ?  ?  ?  :  ?  :  0;  // preset
  ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
  *  0  b  ?  ?  :  1  :  1;  // reduce clear pessimism
  *  0  x  0  ?  :  1  :  1;  // reduce clear pessimism
  0  *  b  ?  ?  :  0  :  0;  // reduce preset pessimism
  0  *  x  1  ?  :  0  :  0;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_IQN_LATCH_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N : QN : QN 
  ?  ?  0  *  ?  :  ?  :  -;  // No change CK=0
  ?  0  1  0  ?  :  ?  :  1;  // Latch 0
  ?  0  *  0  ?  :  1  :  1;  // reduce pessimism when D=0
  1  ?  ?  ?  ?  :  ?  :  1;  // Clear : C dominate P
  0  ?  1  1  ?  :  ?  :  0;  // Latch 1
  0  ?  *  1  ?  :  0  :  0;  // reduce pessimism when D=1
  0  1  ?  ?  ?  :  ?  :  0;  // Preset
  *  0  0  ?  ?  :  1  :  1;   // reduce clear pessimism
  *  0  ?  0  ?  :  1  :  1;   // reduce clear pessimism
  0  *  0  ?  ?  :  0  :  0;   // reduce preset pessimism
  0  *  ?  1  ?  :  0  :  0;   // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;   // notifier
                  
endtable
endprimitive

primitive MGM_L_IQ_FF_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  Q  :  Q 
  ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  0;  // CK in 0
  ?  0  p  0  ?  :  0  :  0;  // reduce pessimism D=0
  1  ?  ?  ?  ?  :  ?  :  0;  // clear: C dominate P
  0  ?  r  1  ?  :  ?  :  1;  // CK in 1
  0  ?  p  1  ?  :  1  :  1;  // reduce pessimism D=1
  0  1  ?  ?  ?  :  ?  :  1;  // preset
  ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
  *  0  b  ?  ?  :  0  :  0;  // reduce clear pessimism
  *  0  x  0  ?  :  0  :  0;  // reduce clear pessimism
  0  *  b  ?  ?  :  1  :  1;  // reduce preset pessimism
  0  *  x  1  ?  :  1  :  1;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_L_IQN_FF_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  QN  :  QN 
  ?  ?  n  ?  ?  :  ?  :  -; // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  1; // CK in 0
  ?  0  p  0  ?  :  1  :  1; // reduce pessimism D=0
  1  0  ?  ?  ?  :  ?  :  1; // clear
  0  ?  r  1  ?  :  ?  :  0; // CK in 1
  0  ?  p  1  ?  :  0  :  0; // reduce pessimism D=1
  ?  1  ?  ?  ?  :  ?  :  0; // preset P dominate C
  ?  ?  b  *  ?  :  ?  :  -; // ignore D change on steady CK : add
  *  0  b  ?  ?  :  1  :  1;  // reduce clear pessimism
  *  0  x  0  ?  :  1  :  1;  // reduce clear pessimism
  0  *  b  ?  ?  :  0  :  0;  // reduce preset pessimism
  0  *  x  1  ?  :  0  :  0;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x; // notifier change
                  
endtable
endprimitive

primitive MGM_L_IQN_LATCH_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N : QN : QN 
  ?  ?  0  *  ?  :  ?  :  -;  // No change CK=0
  ?  0  1  0  ?  :  ?  :  1;  // Latch 0
  ?  0  *  0  ?  :  1  :  1;  // reduce pessimism when D=0
  1  0  ?  ?  ?  :  ?  :  1;  // clear
  0  ?  1  1  ?  :  ?  :  0;  // Latch 1
  0  ?  *  1  ?  :  0  :  0;  // reduce pessimism when D=1
  ?  1  ?  ?  ?  :  ?  :  0;  // Preset P dominate C
  *  0  0  ?  ?  :  1  :  1;   // reduce clear pessimism
  *  0  ?  0  ?  :  1  :  1;   // reduce clear pessimism
  0  *  0  ?  ?  :  0  :  0;   // reduce preset pessimism
  0  *  ?  1  ?  :  0  :  0;   // reduce preset pessimism

//  ?  ?  ?  ?  *  :  ?  :  x;  // notifier
                  
endtable
endprimitive

primitive MOAI22M1HM_udp_0(Z,A1, A2, B1, B2);
  output Z;
  input A1, A2, B1, B2;
  table
  //A1, A2, B1, B2: Z
    0  0  ?  ?: 1;
    ?  ?  1  1: 1;
    1  ?  0  ?: 0;
    1  ?  ?  0: 0;
    ?  1  0  ?: 0;
    ?  1  ?  0: 0;
  endtable
endprimitive

primitive MUX3M0HM_udp_0(Z,A, S0, S1, B, C);
  output Z;
  input A, S0, S1, B, C;
  table
  //A, S0, S1, B, C: Z
    1  0  0  ?  ?: 1;
    ?  1  0  1  ?: 1;
    ?  ?  1  ?  1: 1;
    0  0  0  ?  ?: 0;
    ?  1  0  0  ?: 0;
    ?  ?  1  ?  0: 0;
    1  ?  0  1  ?: 1;
    ?  1  ?  1  1: 1;
    1  0  ?  ?  1: 1;
    1  ?  ?  1  1: 1;
    0  ?  0  0  ?: 0;
    ?  1  ?  0  0: 0;
    0  0  ?  ?  0: 0;
    0  ?  ?  0  0: 0;
  endtable
endprimitive

primitive MUX4M0HM_udp_0(Z,A, S0, S1, B, C, D);
  output Z;
  input A, S0, S1, B, C, D;
  table
  //A, S0, S1, B, C, D: Z
    1  0  0  ?  ?  ?: 1;
    ?  1  0  1  ?  ?: 1;
    ?  0  1  ?  1  ?: 1;
    ?  1  1  ?  ?  1: 1;
    0  0  0  ?  ?  ?: 0;
    ?  1  0  0  ?  ?: 0;
    ?  0  1  ?  0  ?: 0;
    ?  1  1  ?  ?  0: 0;
    1  ?  0  1  ?  ?: 1;
    ?  ?  1  ?  1  1: 1;
    1  0  ?  ?  1  ?: 1;
    ?  1  ?  1  ?  1: 1;
    1  ?  ?  1  1  1: 1;
    0  ?  0  0  ?  ?: 0;
    ?  ?  1  ?  0  0: 0;
    0  0  ?  ?  0  ?: 0;
    ?  1  ?  0  ?  0: 0;
    0  ?  ?  0  0  0: 0;
  endtable
endprimitive

primitive MXB2M0HM_udp_0(Z,A, S, B);
  output Z;
  input A, S, B;
  table
  //A, S, B: Z
    0  0  ?: 1;
    ?  1  0: 1;
    1  0  ?: 0;
    ?  1  1: 0;
    1  ?  1: 0;
    0  ?  0: 1;
  endtable
endprimitive

primitive MXB3M0HM_udp_0(Z,A, S0, S1, B, C);
  output Z;
  input A, S0, S1, B, C;
  table
  //A, S0, S1, B, C: Z
    0  0  0  ?  ?: 1;
    ?  1  0  0  ?: 1;
    ?  ?  1  ?  0: 1;
    1  0  0  ?  ?: 0;
    ?  1  0  1  ?: 0;
    ?  ?  1  ?  1: 0;
    1  ?  0  1  ?: 0;
    ?  1  ?  1  1: 0;
    1  0  ?  ?  1: 0;
    1  ?  ?  1  1: 0;
    0  ?  0  0  ?: 1;
    ?  1  ?  0  0: 1;
    0  0  ?  ?  0: 1;
    0  ?  ?  0  0: 1;
  endtable
endprimitive

primitive MXB4M0HM_udp_0(Z,A, S0, S1, B, C, D);
  output Z;
  input A, S0, S1, B, C, D;
  table
  //A, S0, S1, B, C, D: Z
    0  0  0  ?  ?  ?: 1;
    ?  1  0  0  ?  ?: 1;
    ?  0  1  ?  0  ?: 1;
    ?  1  1  ?  ?  0: 1;
    1  0  0  ?  ?  ?: 0;
    ?  1  0  1  ?  ?: 0;
    ?  0  1  ?  1  ?: 0;
    ?  1  1  ?  ?  1: 0;
    1  ?  0  1  ?  ?: 0;
    ?  ?  1  ?  1  1: 0;
    1  0  ?  ?  1  ?: 0;
    ?  1  ?  1  ?  1: 0;
    1  ?  ?  1  1  1: 0;
    0  ?  0  0  ?  ?: 1;
    ?  ?  1  ?  0  0: 1;
    0  0  ?  ?  0  ?: 1;
    ?  1  ?  0  ?  0: 1;
    0  ?  ?  0  0  0: 1;
  endtable
endprimitive

primitive ND2B1M0HM_udp_0(Z,B, NA);
  output Z;
  input B, NA;
  table
  //B, NA: Z
    0  ?: 1;
    ?  1: 1;
    1  0: 0;
  endtable
endprimitive

primitive ND3B1M0HM_udp_0(Z,B, C, NA);
  output Z;
  input B, C, NA;
  table
  //B, C, NA: Z
    0  ?  ?: 1;
    ?  0  ?: 1;
    ?  ?  1: 1;
    1  1  0: 0;
  endtable
endprimitive

primitive ND3M0HM_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    0  ?  ?: 1;
    ?  0  ?: 1;
    ?  ?  0: 1;
    1  1  1: 0;
  endtable
endprimitive

primitive ND4B1M0HM_udp_0(Z,B, C, D, NA);
  output Z;
  input B, C, D, NA;
  table
  //B, C, D, NA: Z
    0  ?  ?  ?: 1;
    ?  0  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  1: 1;
    1  1  1  0: 0;
  endtable
endprimitive

primitive ND4B2M0HM_udp_0(Z,C, D, NA, NB);
  output Z;
  input C, D, NA, NB;
  table
  //C, D, NA, NB: Z
    0  ?  ?  ?: 1;
    ?  0  ?  ?: 1;
    ?  ?  1  ?: 1;
    ?  ?  ?  1: 1;
    1  1  0  0: 0;
  endtable
endprimitive

primitive ND4M0HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    0  ?  ?  ?: 1;
    ?  0  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  0: 1;
    1  1  1  1: 0;
  endtable
endprimitive

primitive NR2B1M0HM_udp_0(Z,B, NA);
  output Z;
  input B, NA;
  table
  //B, NA: Z
    0  1: 1;
    1  ?: 0;
    ?  0: 0;
  endtable
endprimitive

primitive NR3B1M0HM_udp_0(Z,B, C, NA);
  output Z;
  input B, C, NA;
  table
  //B, C, NA: Z
    0  0  1: 1;
    1  ?  ?: 0;
    ?  1  ?: 0;
    ?  ?  0: 0;
  endtable
endprimitive

primitive NR3M0HM_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    0  0  0: 1;
    1  ?  ?: 0;
    ?  1  ?: 0;
    ?  ?  1: 0;
  endtable
endprimitive

primitive NR4B1M0HM_udp_0(Z,B, C, D, NA);
  output Z;
  input B, C, D, NA;
  table
  //B, C, D, NA: Z
    0  0  0  1: 1;
    1  ?  ?  ?: 0;
    ?  1  ?  ?: 0;
    ?  ?  1  ?: 0;
    ?  ?  ?  0: 0;
  endtable
endprimitive

primitive NR4B2M0HM_udp_0(Z,C, D, NA, NB);
  output Z;
  input C, D, NA, NB;
  table
  //C, D, NA, NB: Z
    0  0  1  1: 1;
    1  ?  ?  ?: 0;
    ?  1  ?  ?: 0;
    ?  ?  0  ?: 0;
    ?  ?  ?  0: 0;
  endtable
endprimitive

primitive NR4M0HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    0  0  0  0: 1;
    1  ?  ?  ?: 0;
    ?  1  ?  ?: 0;
    ?  ?  1  ?: 0;
    ?  ?  ?  1: 0;
  endtable
endprimitive

primitive OA211M12HM_udp_0(Z,A1, B, C, A2);
  output Z;
  input A1, B, C, A2;
  table
  //A1, B, C, A2: Z
    1  1  1  ?: 1;
    ?  1  1  1: 1;
    0  ?  ?  0: 0;
    ?  0  ?  ?: 0;
    ?  ?  0  ?: 0;
  endtable
endprimitive

primitive OA21M0HM_udp_0(Z,A1, B, A2);
  output Z;
  input A1, B, A2;
  table
  //A1, B, A2: Z
    1  1  ?: 1;
    ?  1  1: 1;
    0  ?  0: 0;
    ?  0  ?: 0;
  endtable
endprimitive

primitive OA221M1HM_udp_0(Z,A1, B1, C, B2, A2);
  output Z;
  input A1, B1, C, B2, A2;
  table
  //A1, B1, C, B2, A2: Z
    1  1  1  ?  ?: 1;
    1  ?  1  1  ?: 1;
    ?  1  1  ?  1: 1;
    ?  ?  1  1  1: 1;
    0  ?  ?  ?  0: 0;
    ?  0  ?  0  ?: 0;
    ?  ?  0  ?  ?: 0;
  endtable
endprimitive

primitive OA222M1HM_udp_0(Z,A1, B1, C1, C2, B2, A2);
  output Z;
  input A1, B1, C1, C2, B2, A2;
  table
  //A1, B1, C1, C2, B2, A2: Z
    1  1  1  ?  ?  ?: 1;
    1  1  ?  1  ?  ?: 1;
    1  ?  1  ?  1  ?: 1;
    1  ?  ?  1  1  ?: 1;
    ?  1  1  ?  ?  1: 1;
    ?  1  ?  1  ?  1: 1;
    ?  ?  1  ?  1  1: 1;
    ?  ?  ?  1  1  1: 1;
    0  ?  ?  ?  ?  0: 0;
    ?  0  ?  ?  0  ?: 0;
    ?  ?  0  0  ?  ?: 0;
  endtable
endprimitive

primitive OA22M0HM_udp_0(Z,A1, B1, B2, A2);
  output Z;
  input A1, B1, B2, A2;
  table
  //A1, B1, B2, A2: Z
    1  1  ?  ?: 1;
    1  ?  1  ?: 1;
    ?  1  ?  1: 1;
    ?  ?  1  1: 1;
    0  ?  ?  0: 0;
    ?  0  0  ?: 0;
  endtable
endprimitive

primitive OA31M1HM_udp_0(Z,A1, B, A2, A3);
  output Z;
  input A1, B, A2, A3;
  table
  //A1, B, A2, A3: Z
    1  1  ?  ?: 1;
    ?  1  1  ?: 1;
    ?  1  ?  1: 1;
    0  ?  0  0: 0;
    ?  0  ?  ?: 0;
  endtable
endprimitive

primitive OA32M1HM_udp_0(Z,A1, B1, B2, A2, A3);
  output Z;
  input A1, B1, B2, A2, A3;
  table
  //A1, B1, B2, A2, A3: Z
    1  1  ?  ?  ?: 1;
    1  ?  1  ?  ?: 1;
    ?  1  ?  1  ?: 1;
    ?  ?  1  1  ?: 1;
    ?  1  ?  ?  1: 1;
    ?  ?  1  ?  1: 1;
    0  ?  ?  0  0: 0;
    ?  0  0  ?  ?: 0;
  endtable
endprimitive

primitive OA33M1HM_udp_0(Z,A1, B1, B2, B3, A2, A3);
  output Z;
  input A1, B1, B2, B3, A2, A3;
  table
  //A1, B1, B2, B3, A2, A3: Z
    1  1  ?  ?  ?  ?: 1;
    1  ?  1  ?  ?  ?: 1;
    1  ?  ?  1  ?  ?: 1;
    ?  1  ?  ?  1  ?: 1;
    ?  ?  1  ?  1  ?: 1;
    ?  ?  ?  1  1  ?: 1;
    ?  1  ?  ?  ?  1: 1;
    ?  ?  1  ?  ?  1: 1;
    ?  ?  ?  1  ?  1: 1;
    0  ?  ?  ?  0  0: 0;
    ?  0  0  0  ?  ?: 0;
  endtable
endprimitive

primitive OAI211B100M0HM_udp_0(Z,A1, NA2, B, C);
  output Z;
  input A1, NA2, B, C;
  table
  //A1, NA2, B, C: Z
    0  1  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  0: 1;
    1  ?  1  1: 0;
    ?  0  1  1: 0;
  endtable
endprimitive

primitive OAI211M0HM_udp_0(Z,A1, A2, B, C);
  output Z;
  input A1, A2, B, C;
  table
  //A1, A2, B, C: Z
    0  0  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  0: 1;
    1  ?  1  1: 0;
    ?  1  1  1: 0;
  endtable
endprimitive

primitive OAI21B10M0HM_udp_0(Z,A1, NA2, B);
  output Z;
  input A1, NA2, B;
  table
  //A1, NA2, B: Z
    0  1  ?: 1;
    ?  ?  0: 1;
    1  ?  1: 0;
    ?  0  1: 0;
  endtable
endprimitive

primitive OAI21B20M0HM_udp_0(Z,B, NA1, NA2);
  output Z;
  input B, NA1, NA2;
  table
  //B, NA1, NA2: Z
    0  ?  ?: 1;
    ?  1  1: 1;
    1  0  ?: 0;
    1  ?  0: 0;
  endtable
endprimitive

primitive OAI21M0HM_udp_0(Z,A1, A2, B);
  output Z;
  input A1, A2, B;
  table
  //A1, A2, B: Z
    0  0  ?: 1;
    ?  ?  0: 1;
    1  ?  1: 0;
    ?  1  1: 0;
  endtable
endprimitive

primitive OAI221M0HM_udp_0(Z,A1, A2, B1, B2, C);
  output Z;
  input A1, A2, B1, B2, C;
  table
  //A1, A2, B1, B2, C: Z
    0  0  ?  ?  ?: 1;
    ?  ?  0  0  ?: 1;
    ?  ?  ?  ?  0: 1;
    1  ?  1  ?  1: 0;
    1  ?  ?  1  1: 0;
    ?  1  1  ?  1: 0;
    ?  1  ?  1  1: 0;
  endtable
endprimitive

primitive OAI222M0HM_udp_0(Z,A1, A2, B1, B2, C1, C2);
  output Z;
  input A1, A2, B1, B2, C1, C2;
  table
  //A1, A2, B1, B2, C1, C2: Z
    0  0  ?  ?  ?  ?: 1;
    ?  ?  0  0  ?  ?: 1;
    ?  ?  ?  ?  0  0: 1;
    1  ?  1  ?  1  ?: 0;
    1  ?  1  ?  ?  1: 0;
    1  ?  ?  1  1  ?: 0;
    1  ?  ?  1  ?  1: 0;
    ?  1  1  ?  1  ?: 0;
    ?  1  1  ?  ?  1: 0;
    ?  1  ?  1  1  ?: 0;
    ?  1  ?  1  ?  1: 0;
  endtable
endprimitive

primitive OAI22B10M0HM_udp_0(Z,A1, NA2, B1, B2);
  output Z;
  input A1, NA2, B1, B2;
  table
  //A1, NA2, B1, B2: Z
    0  1  ?  ?: 1;
    ?  ?  0  0: 1;
    1  ?  1  ?: 0;
    1  ?  ?  1: 0;
    ?  0  1  ?: 0;
    ?  0  ?  1: 0;
  endtable
endprimitive

primitive OAI22M0HM_udp_0(Z,A1, A2, B1, B2);
  output Z;
  input A1, A2, B1, B2;
  table
  //A1, A2, B1, B2: Z
    0  0  ?  ?: 1;
    ?  ?  0  0: 1;
    1  ?  1  ?: 0;
    1  ?  ?  1: 0;
    ?  1  1  ?: 0;
    ?  1  ?  1: 0;
  endtable
endprimitive

primitive OAI31M0HM_udp_0(Z,A1, A2, A3, B);
  output Z;
  input A1, A2, A3, B;
  table
  //A1, A2, A3, B: Z
    0  0  0  ?: 1;
    ?  ?  ?  0: 1;
    1  ?  ?  1: 0;
    ?  1  ?  1: 0;
    ?  ?  1  1: 0;
  endtable
endprimitive

primitive OAI32M0HM_udp_0(Z,A1, A2, A3, B1, B2);
  output Z;
  input A1, A2, A3, B1, B2;
  table
  //A1, A2, A3, B1, B2: Z
    0  0  0  ?  ?: 1;
    ?  ?  ?  0  0: 1;
    1  ?  ?  1  ?: 0;
    1  ?  ?  ?  1: 0;
    ?  1  ?  1  ?: 0;
    ?  1  ?  ?  1: 0;
    ?  ?  1  1  ?: 0;
    ?  ?  1  ?  1: 0;
  endtable
endprimitive

primitive OAI33M0HM_udp_0(Z,A1, A2, A3, B1, B2, B3);
  output Z;
  input A1, A2, A3, B1, B2, B3;
  table
  //A1, A2, A3, B1, B2, B3: Z
    0  0  0  ?  ?  ?: 1;
    ?  ?  ?  0  0  0: 1;
    1  ?  ?  1  ?  ?: 0;
    1  ?  ?  ?  1  ?: 0;
    1  ?  ?  ?  ?  1: 0;
    ?  1  ?  1  ?  ?: 0;
    ?  1  ?  ?  1  ?: 0;
    ?  1  ?  ?  ?  1: 0;
    ?  ?  1  1  ?  ?: 0;
    ?  ?  1  ?  1  ?: 0;
    ?  ?  1  ?  ?  1: 0;
  endtable
endprimitive

primitive OR2M0HM_udp_0(Z,A, B);
  output Z;
  input A, B;
  table
  //A, B: Z
    1  ?: 1;
    ?  1: 1;
    0  0: 0;
  endtable
endprimitive

primitive OR3M0HM_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    1  ?  ?: 1;
    ?  1  ?: 1;
    ?  ?  1: 1;
    0  0  0: 0;
  endtable
endprimitive

primitive OR4M0HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  ?  ?  ?: 1;
    ?  1  ?  ?: 1;
    ?  ?  1  ?: 1;
    ?  ?  ?  1: 1;
    0  0  0  0: 0;
  endtable
endprimitive

primitive OR6M12HM_udp_0(Z,A, B, C, D, E, F);
  output Z;
  input A, B, C, D, E, F;
  table
  //A, B, C, D, E, F: Z
    1  ?  ?  ?  ?  ?: 1;
    ?  1  ?  ?  ?  ?: 1;
    ?  ?  1  ?  ?  ?: 1;
    ?  ?  ?  1  ?  ?: 1;
    ?  ?  ?  ?  1  ?: 1;
    ?  ?  ?  ?  ?  1: 1;
    0  0  0  0  0  0: 0;
  endtable
endprimitive

primitive SDFAQM1HM_udp_0(MGM_D,A, B, SE, SD);
  output MGM_D;
  input A, B, SE, SD;
  table
  //A, B, SE, SD: MGM_D
    1  1  0  ?: 1;
    ?  ?  1  1: 1;
    0  ?  0  ?: 0;
    ?  0  0  ?: 0;
    ?  ?  1  0: 0;
    1  1  ?  1: 1;
    0  ?  ?  0: 0;
    ?  0  ?  0: 0;
  endtable
endprimitive

primitive SDFEM1HM_udp_0(MGM_D,D, E, SE, IQ, SD);
  output MGM_D;
  input D, E, SE, IQ, SD;
  table
  //D, E, SE, IQ, SD: MGM_D
    1  1  0  ?  ?: 1;
    1  ?  0  1  ?: 1;
    ?  0  0  1  ?: 1;
    ?  ?  1  ?  1: 1;
    0  1  0  ?  ?: 0;
    0  ?  0  0  ?: 0;
    ?  0  0  0  ?: 0;
    ?  ?  1  ?  0: 0;
    1  1  ?  ?  1: 1;
    1  ?  ?  1  1: 1;
    ?  0  ?  1  1: 1;
    0  1  ?  ?  0: 0;
    0  ?  ?  0  0: 0;
    ?  0  ?  0  0: 0;
  endtable
endprimitive

primitive SDFEQZRM1HM_udp_0(MGM_D,D, E, RB, SE, IQ, SD);
  output MGM_D;
  input D, E, RB, SE, IQ, SD;
  table
  //D, E, RB, SE, IQ, SD: MGM_D
    1  1  1  0  ?  ?: 1;
    1  ?  1  0  1  ?: 1;
    ?  0  1  0  1  ?: 1;
    ?  ?  ?  1  ?  1: 1;
    0  1  ?  0  ?  ?: 0;
    0  ?  ?  0  0  ?: 0;
    ?  0  ?  0  0  ?: 0;
    ?  ?  0  0  ?  ?: 0;
    ?  ?  ?  1  ?  0: 0;
    1  1  1  ?  ?  1: 1;
    1  ?  1  ?  1  1: 1;
    ?  0  1  ?  1  1: 1;
    0  1  ?  ?  ?  0: 0;
    0  ?  ?  ?  0  0: 0;
    ?  0  ?  ?  0  0: 0;
    ?  ?  0  ?  ?  0: 0;
  endtable
endprimitive

primitive SDFMM1HM_udp_0(MGM_D,D1, S, SE, D2, SD);
  output MGM_D;
  input D1, S, SE, D2, SD;
  table
  //D1, S, SE, D2, SD: MGM_D
    1  1  0  ?  ?: 1;
    ?  0  0  1  ?: 1;
    ?  ?  1  ?  1: 1;
    0  1  0  ?  ?: 0;
    ?  0  0  0  ?: 0;
    ?  ?  1  ?  0: 0;
    1  1  ?  ?  1: 1;
    ?  0  ?  1  1: 1;
    0  1  ?  ?  0: 0;
    ?  0  ?  0  0: 0;
    1  ?  0  1  ?: 1;
    0  ?  0  0  ?: 0;
    1  ?  ?  1  1: 1;
    0  ?  ?  0  0: 0;
  endtable
endprimitive

primitive XNR4M1HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  1  1  1: 1;
    1  1  0  0: 1;
    1  0  1  0: 1;
    1  0  0  1: 1;
    0  1  1  0: 1;
    0  1  0  1: 1;
    0  0  1  1: 1;
    0  0  0  0: 1;
    1  1  1  0: 0;
    1  1  0  1: 0;
    1  0  1  1: 0;
    1  0  0  0: 0;
    0  1  1  1: 0;
    0  1  0  0: 0;
    0  0  1  0: 0;
    0  0  0  1: 0;
  endtable
endprimitive

primitive XOR4M1HM_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  1  1  0: 1;
    1  1  0  1: 1;
    1  0  1  1: 1;
    1  0  0  0: 1;
    0  1  1  1: 1;
    0  1  0  0: 1;
    0  0  1  0: 1;
    0  0  0  1: 1;
    1  1  1  1: 0;
    1  1  0  0: 0;
    1  0  1  0: 0;
    1  0  0  1: 0;
    0  1  1  0: 0;
    0  1  0  1: 0;
    0  0  1  1: 0;
    0  0  0  0: 0;
  endtable
endprimitive
